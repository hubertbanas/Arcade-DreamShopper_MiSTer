library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"F0",X"4F",X"E7",X"C3",X"B4",X"01",X"FF",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"FF",X"FF",
		X"D5",X"07",X"5F",X"16",X"00",X"19",X"D1",X"C9",X"E1",X"18",X"33",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"AF",X"32",X"00",X"50",X"32",X"C0",X"50",X"C9",X"E7",X"3E",X"01",X"32",X"00",X"50",X"C9",X"FF",
		X"18",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CD",X"AA",X"01",X"0F",X"0F",X"0F",X"E6",X"1E",
		X"5F",X"16",X"00",X"21",X"D4",X"01",X"19",X"5E",X"23",X"56",X"EB",X"F1",X"F5",X"E9",X"CB",X"27",
		X"5F",X"16",X"00",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"ED",X"73",X"1C",X"48",X"31",X"90",X"4F",X"08",X"D9",X"E7",
		X"DD",X"E5",X"FD",X"E5",X"CD",X"E8",X"01",X"FD",X"E1",X"DD",X"E1",X"0E",X"03",X"21",X"B0",X"4B",
		X"06",X"09",X"11",X"06",X"00",X"7E",X"FE",X"01",X"23",X"20",X"1B",X"79",X"A6",X"23",X"28",X"03",
		X"35",X"28",X"0C",X"19",X"10",X"EF",X"EF",X"D9",X"08",X"ED",X"7B",X"1C",X"48",X"ED",X"45",X"2B",
		X"CB",X"FE",X"2B",X"36",X"03",X"23",X"23",X"18",X"EA",X"31",X"F0",X"4F",X"FB",X"0E",X"00",X"21",
		X"B0",X"4B",X"06",X"09",X"11",X"08",X"00",X"7E",X"CB",X"7F",X"20",X"04",X"FE",X"02",X"30",X"06",
		X"0C",X"19",X"10",X"F3",X"18",X"E7",X"F3",X"79",X"32",X"00",X"48",X"7E",X"36",X"02",X"23",X"CB",
		X"BE",X"23",X"36",X"00",X"23",X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"23",X"EB",X"FE",X"04",
		X"20",X"04",X"50",X"59",X"FB",X"E9",X"F9",X"FE",X"02",X"28",X"04",X"1A",X"C1",X"18",X"01",X"F1",
		X"C1",X"D1",X"E1",X"FD",X"E1",X"DD",X"E1",X"FB",X"C9",X"CD",X"9A",X"01",X"36",X"04",X"23",X"72",
		X"23",X"72",X"23",X"71",X"23",X"70",X"18",X"E7",X"CD",X"9A",X"01",X"72",X"18",X"E1",X"CD",X"97",
		X"01",X"7E",X"FE",X"02",X"C2",X"A9",X"00",X"23",X"7E",X"CB",X"7F",X"20",X"15",X"E6",X"40",X"4F",
		X"F1",X"F5",X"E6",X"0F",X"B1",X"77",X"23",X"70",X"2B",X"2B",X"36",X"01",X"CD",X"89",X"01",X"C3",
		X"A9",X"00",X"CB",X"BE",X"1E",X"06",X"19",X"7E",X"18",X"B2",X"CD",X"9A",X"01",X"CB",X"BE",X"7E",
		X"B7",X"28",X"AC",X"FE",X"04",X"28",X"A8",X"1E",X"07",X"19",X"70",X"11",X"FA",X"FF",X"19",X"CB",
		X"F6",X"CB",X"FE",X"FE",X"01",X"20",X"98",X"2B",X"36",X"03",X"18",X"93",X"CD",X"9A",X"01",X"7E",
		X"B7",X"28",X"8C",X"CB",X"FE",X"18",X"88",X"CD",X"97",X"01",X"72",X"C3",X"A9",X"00",X"CD",X"9A",
		X"01",X"1E",X"05",X"19",X"71",X"23",X"70",X"C3",X"EF",X"00",X"CD",X"97",X"01",X"23",X"CB",X"76",
		X"CB",X"B6",X"1E",X"06",X"19",X"7E",X"C3",X"EC",X"00",X"01",X"03",X"00",X"09",X"EB",X"21",X"02",
		X"00",X"39",X"EB",X"73",X"23",X"72",X"C9",X"3A",X"00",X"48",X"E6",X"0F",X"21",X"B0",X"4B",X"16",
		X"00",X"5F",X"CB",X"23",X"CB",X"23",X"CB",X"23",X"19",X"C9",X"DD",X"E3",X"FD",X"E5",X"E5",X"D5",
		X"C5",X"F5",X"DD",X"E9",X"21",X"00",X"40",X"01",X"00",X"20",X"36",X"00",X"23",X"0B",X"78",X"B1",
		X"20",X"F8",X"3A",X"00",X"50",X"2F",X"CB",X"7F",X"C2",X"00",X"A7",X"3E",X"00",X"01",X"F0",X"2E",
		X"FF",X"C3",X"A9",X"00",X"F9",X"00",X"08",X"01",X"0E",X"01",X"0E",X"01",X"3A",X"01",X"5C",X"01",
		X"67",X"01",X"6E",X"01",X"7A",X"01",X"FF",X"FF",X"3A",X"02",X"48",X"CB",X"67",X"C0",X"3A",X"C0",
		X"50",X"2F",X"32",X"1A",X"48",X"21",X"80",X"50",X"36",X"01",X"36",X"00",X"21",X"1E",X"48",X"7E",
		X"CB",X"BF",X"B7",X"28",X"0B",X"3D",X"CB",X"FF",X"77",X"20",X"05",X"AF",X"77",X"32",X"07",X"50",
		X"3A",X"00",X"50",X"2F",X"E6",X"A0",X"57",X"21",X"03",X"48",X"7E",X"B7",X"7A",X"16",X"A0",X"20",
		X"1C",X"A2",X"CA",X"BD",X"02",X"FE",X"20",X"20",X"07",X"E5",X"21",X"1E",X"48",X"CB",X"FE",X"E1",
		X"36",X"24",X"C3",X"BD",X"02",X"00",X"00",X"00",X"01",X"00",X"02",X"00",X"03",X"35",X"28",X"14",
		X"4F",X"7E",X"FE",X"22",X"79",X"30",X"06",X"A2",X"C2",X"BD",X"02",X"18",X"0B",X"A2",X"C2",X"BD",
		X"02",X"C3",X"00",X"00",X"A2",X"C2",X"00",X"00",X"36",X"00",X"3A",X"1E",X"48",X"CB",X"7F",X"28",
		X"0A",X"3E",X"06",X"32",X"1E",X"48",X"3E",X"01",X"32",X"07",X"50",X"06",X"64",X"21",X"04",X"48",
		X"4E",X"23",X"7E",X"81",X"B8",X"30",X"13",X"06",X"00",X"77",X"21",X"36",X"02",X"CB",X"21",X"09",
		X"11",X"07",X"48",X"06",X"02",X"CD",X"DA",X"8F",X"18",X"08",X"05",X"70",X"21",X"09",X"09",X"22",
		X"06",X"48",X"3A",X"02",X"48",X"CB",X"7F",X"20",X"15",X"3E",X"0E",X"CD",X"40",X"03",X"21",X"49",
		X"42",X"DD",X"21",X"06",X"48",X"1E",X"02",X"06",X"02",X"0E",X"FF",X"CD",X"1E",X"90",X"21",X"01",
		X"48",X"CB",X"7E",X"CB",X"FE",X"20",X"06",X"3E",X"00",X"01",X"F2",X"2E",X"FF",X"21",X"40",X"48",
		X"DD",X"21",X"F0",X"4F",X"FD",X"21",X"60",X"50",X"06",X"08",X"CB",X"7E",X"20",X"4F",X"4E",X"0C",
		X"3A",X"1B",X"48",X"57",X"CB",X"FE",X"23",X"7E",X"CB",X"42",X"28",X"09",X"EE",X"C0",X"E6",X"C0",
		X"5F",X"3E",X"3F",X"A6",X"B3",X"07",X"07",X"DD",X"77",X"00",X"23",X"7E",X"CB",X"42",X"28",X"04",
		X"ED",X"44",X"C6",X"10",X"D6",X"02",X"FD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",X"23",X"7E",
		X"CB",X"42",X"28",X"04",X"ED",X"44",X"C6",X"10",X"FD",X"77",X"01",X"23",X"DD",X"23",X"DD",X"23",
		X"FD",X"23",X"FD",X"23",X"05",X"CA",X"68",X"03",X"0D",X"28",X"AF",X"18",X"B3",X"11",X"05",X"00",
		X"19",X"DD",X"23",X"DD",X"23",X"FD",X"23",X"FD",X"23",X"10",X"9F",X"C3",X"68",X"03",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"47",X"00",X"00",X"00",X"FE",X"0E",X"20",X"09",X"3A",X"02",X"48",X"CB",X"7F",X"78",X"C0",X"18",
		X"07",X"3A",X"01",X"48",X"CB",X"7F",X"78",X"C8",X"D5",X"E5",X"DD",X"E5",X"FD",X"E5",X"CD",X"6E",
		X"04",X"FD",X"E1",X"DD",X"E1",X"E1",X"D1",X"C9",X"C3",X"6B",X"03",X"DD",X"21",X"20",X"48",X"DD",
		X"E5",X"FD",X"E1",X"DD",X"23",X"DD",X"23",X"0E",X"03",X"06",X"01",X"DD",X"CB",X"00",X"7E",X"C5",
		X"DD",X"E5",X"C4",X"93",X"03",X"DD",X"E1",X"C1",X"11",X"0A",X"00",X"DD",X"19",X"CB",X"20",X"0D",
		X"20",X"E9",X"C9",X"DD",X"35",X"07",X"C0",X"DD",X"7E",X"02",X"DD",X"77",X"07",X"DD",X"CB",X"00",
		X"46",X"28",X"08",X"DD",X"35",X"08",X"C0",X"DD",X"CB",X"00",X"86",X"DD",X"CB",X"00",X"4E",X"28",
		X"08",X"DD",X"35",X"08",X"C0",X"DD",X"CB",X"00",X"8E",X"DD",X"6E",X"05",X"DD",X"66",X"06",X"7E",
		X"23",X"DD",X"75",X"05",X"DD",X"74",X"06",X"CB",X"7F",X"20",X"07",X"DD",X"77",X"09",X"CD",X"CC",
		X"05",X"C9",X"FE",X"80",X"20",X"01",X"C9",X"FE",X"C0",X"20",X"0D",X"4E",X"23",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"CD",X"3A",X"05",X"18",X"D1",X"FE",X"C1",X"20",X"05",X"CD",X"4B",X"05",X"18",
		X"C8",X"4F",X"E6",X"F0",X"FE",X"A0",X"20",X"05",X"CD",X"88",X"05",X"18",X"BC",X"FE",X"90",X"20",
		X"05",X"CD",X"75",X"05",X"18",X"B3",X"FE",X"E0",X"20",X"0C",X"EB",X"CD",X"55",X"05",X"DD",X"73",
		X"05",X"DD",X"72",X"06",X"18",X"A3",X"FE",X"D0",X"20",X"0E",X"79",X"E6",X"0F",X"DD",X"77",X"08",
		X"DD",X"CB",X"00",X"C6",X"CD",X"A2",X"05",X"C9",X"FE",X"B0",X"20",X"0B",X"79",X"E6",X"0F",X"DD",
		X"77",X"08",X"DD",X"CB",X"00",X"CE",X"C9",X"FE",X"F0",X"20",X"FC",X"CD",X"FB",X"04",X"DD",X"CB",
		X"00",X"76",X"20",X"09",X"DD",X"E5",X"E1",X"06",X"0A",X"CD",X"C6",X"05",X"C9",X"DD",X"CB",X"00",
		X"FE",X"DD",X"4E",X"02",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"DD",X"71",X"07",X"DD",X"75",X"05",
		X"DD",X"74",X"06",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"C3",X"B9",X"03",X"DD",X"21",
		X"90",X"9C",X"FD",X"21",X"20",X"48",X"CB",X"7F",X"28",X"09",X"E6",X"0F",X"CA",X"D5",X"04",X"47",
		X"C3",X"FB",X"04",X"16",X"00",X"3D",X"CB",X"27",X"5F",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",
		X"01",X"E5",X"DD",X"E1",X"DD",X"7E",X"00",X"E6",X"0E",X"47",X"CD",X"1F",X"06",X"E5",X"06",X"0A",
		X"CD",X"C6",X"05",X"E1",X"CB",X"FE",X"DD",X"CB",X"00",X"76",X"28",X"02",X"CB",X"F6",X"23",X"DD",
		X"7E",X"01",X"77",X"23",X"DD",X"7E",X"02",X"77",X"23",X"DD",X"4E",X"03",X"71",X"23",X"DD",X"46",
		X"04",X"70",X"23",X"71",X"23",X"70",X"23",X"36",X"01",X"DD",X"CB",X"00",X"7E",X"C0",X"01",X"05",
		X"00",X"DD",X"09",X"18",X"BF",X"21",X"20",X"48",X"06",X"20",X"CD",X"C6",X"05",X"01",X"00",X"00",
		X"1E",X"07",X"CD",X"94",X"05",X"04",X"1D",X"20",X"F9",X"0E",X"FF",X"CD",X"94",X"05",X"04",X"0E",
		X"00",X"1E",X"08",X"CD",X"94",X"05",X"04",X"1D",X"20",X"F9",X"C9",X"0E",X"00",X"CD",X"88",X"05",
		X"78",X"FD",X"4E",X"00",X"FE",X"01",X"20",X"06",X"CB",X"81",X"CB",X"99",X"18",X"0E",X"FE",X"02",
		X"20",X"06",X"CB",X"89",X"CB",X"A1",X"18",X"04",X"CB",X"91",X"CB",X"A9",X"21",X"25",X"05",X"E5",
		X"C5",X"79",X"C3",X"BA",X"05",X"C5",X"CB",X"38",X"CB",X"20",X"0E",X"00",X"CD",X"94",X"05",X"04",
		X"CD",X"94",X"05",X"C1",X"CD",X"1F",X"06",X"CB",X"BE",X"C9",X"C5",X"06",X"06",X"CD",X"94",X"05",
		X"C1",X"C5",X"78",X"07",X"07",X"07",X"FD",X"B6",X"00",X"18",X"6F",X"C5",X"78",X"07",X"07",X"07",
		X"FD",X"AE",X"00",X"18",X"65",X"C5",X"06",X"0B",X"1A",X"4F",X"13",X"CD",X"94",X"05",X"04",X"1A",
		X"4F",X"13",X"CD",X"94",X"05",X"C1",X"C5",X"0E",X"10",X"CD",X"88",X"05",X"C1",X"C5",X"06",X"0D",
		X"CD",X"94",X"05",X"C1",X"C9",X"0E",X"00",X"C5",X"06",X"0B",X"CD",X"94",X"05",X"04",X"CD",X"94",
		X"05",X"04",X"CD",X"94",X"05",X"C1",X"18",X"00",X"C5",X"CB",X"38",X"3E",X"08",X"80",X"47",X"CD",
		X"94",X"05",X"C1",X"C9",X"78",X"D3",X"07",X"79",X"D3",X"06",X"C9",X"C5",X"78",X"FD",X"B6",X"00",
		X"18",X"18",X"C5",X"78",X"FD",X"4E",X"00",X"FE",X"01",X"20",X"04",X"CB",X"81",X"18",X"0A",X"FE",
		X"02",X"20",X"04",X"CB",X"89",X"18",X"02",X"CB",X"91",X"79",X"FD",X"77",X"00",X"2F",X"4F",X"06",
		X"07",X"CD",X"94",X"05",X"C1",X"C9",X"AF",X"77",X"23",X"10",X"FC",X"C9",X"4F",X"DD",X"7E",X"01",
		X"B7",X"28",X"18",X"CB",X"7F",X"20",X"0C",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"81",
		X"4F",X"18",X"08",X"5F",X"79",X"C6",X"10",X"1C",X"20",X"FB",X"4F",X"21",X"3B",X"06",X"59",X"CB",
		X"3B",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"CB",X"23",X"16",X"00",X"19",X"5E",X"23",X"56",X"79",
		X"E6",X"0F",X"6F",X"CB",X"25",X"26",X"00",X"19",X"EB",X"C5",X"CB",X"38",X"CB",X"20",X"1A",X"4F",
		X"13",X"CD",X"94",X"05",X"04",X"1A",X"4F",X"CD",X"94",X"05",X"C1",X"CD",X"9B",X"05",X"C9",X"C5",
		X"FD",X"E5",X"D1",X"CB",X"38",X"CB",X"20",X"48",X"06",X"00",X"21",X"35",X"06",X"09",X"4E",X"23",
		X"46",X"EB",X"09",X"C1",X"C9",X"02",X"00",X"0C",X"00",X"16",X"00",X"4B",X"06",X"63",X"06",X"7B",
		X"06",X"93",X"06",X"AB",X"06",X"C3",X"06",X"DB",X"06",X"F3",X"06",X"5D",X"0D",X"9C",X"0C",X"E7",
		X"0B",X"3C",X"0B",X"9B",X"0A",X"02",X"0A",X"73",X"09",X"EB",X"08",X"6B",X"08",X"F2",X"07",X"80",
		X"07",X"14",X"07",X"AE",X"06",X"4E",X"06",X"F4",X"05",X"9E",X"05",X"4D",X"05",X"01",X"05",X"B9",
		X"04",X"75",X"04",X"35",X"04",X"F9",X"03",X"C0",X"03",X"8A",X"03",X"57",X"03",X"27",X"03",X"FA",
		X"02",X"CF",X"02",X"A7",X"02",X"81",X"02",X"5D",X"02",X"3B",X"02",X"1B",X"02",X"FC",X"01",X"E0",
		X"01",X"C5",X"01",X"AC",X"01",X"94",X"01",X"7D",X"01",X"68",X"01",X"53",X"01",X"40",X"01",X"2E",
		X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E2",X"00",X"D6",X"00",X"CA",X"00",X"BE",
		X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",X"00",X"78",
		X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",X"00",X"4C",
		X"00",X"47",X"00",X"43",X"00",X"40",X"00",X"3C",X"00",X"39",X"00",X"35",X"00",X"32",X"00",X"30",
		X"00",X"2D",X"00",X"2A",X"00",X"28",X"00",X"26",X"00",X"24",X"00",X"22",X"00",X"20",X"00",X"1E",
		X"00",X"1C",X"00",X"1B",X"00",X"19",X"00",X"18",X"00",X"16",X"00",X"15",X"00",X"14",X"00",X"13",
		X"00",X"12",X"00",X"11",X"00",X"10",X"00",X"0F",X"00",X"0E",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1C",X"0D",X"A0",X"03",X"A1",X"01",X"A2",X"0B",X"A0",X"1C",X"01",X"A0",X"01",X"A3",X"0B",X"A4",
		X"03",X"A5",X"01",X"AC",X"09",X"A4",X"01",X"A6",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",
		X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",
		X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",
		X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",
		X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",
		X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",
		X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A4",X"01",X"A5",X"98",X"01",X"AC",X"01",X"A4",X"1C",X"9C",
		X"1C",X"9C",X"1C",X"01",X"A7",X"01",X"A8",X"98",X"01",X"A9",X"01",X"A7",X"1C",X"01",X"A0",X"01",
		X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",
		X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",
		X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",
		X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",
		X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",
		X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",
		X"1C",X"01",X"A0",X"01",X"A1",X"98",X"01",X"A2",X"01",X"A0",X"1C",X"01",X"A0",X"01",X"AA",X"0B",
		X"A7",X"03",X"A8",X"01",X"A9",X"09",X"A7",X"01",X"AB",X"01",X"A0",X"1C",X"0D",X"A0",X"03",X"A1",
		X"01",X"A2",X"0B",X"A0",X"00",X"4D",X"08",X"57",X"08",X"6A",X"08",X"74",X"08",X"87",X"08",X"9A",
		X"08",X"AD",X"08",X"BA",X"08",X"CD",X"08",X"E0",X"08",X"FC",X"08",X"09",X"09",X"1C",X"09",X"38",
		X"09",X"4B",X"09",X"58",X"09",X"6B",X"09",X"7E",X"09",X"91",X"09",X"9E",X"09",X"20",X"AA",X"AA",
		X"01",X"FF",X"10",X"01",X"01",X"10",X"FF",X"34",X"AA",X"AA",X"02",X"FE",X"04",X"02",X"FF",X"08",
		X"01",X"00",X"04",X"02",X"01",X"08",X"02",X"02",X"04",X"FF",X"40",X"AA",X"AA",X"02",X"FF",X"10",
		X"02",X"01",X"10",X"FF",X"28",X"AA",X"AA",X"01",X"FE",X"0A",X"01",X"FF",X"05",X"01",X"00",X"02",
		X"01",X"01",X"05",X"01",X"02",X"12",X"FF",X"30",X"AA",X"AA",X"01",X"FE",X"12",X"01",X"FF",X"05",
		X"01",X"00",X"02",X"01",X"01",X"05",X"01",X"02",X"12",X"FF",X"38",X"AA",X"AA",X"01",X"FE",X"12",
		X"01",X"FF",X"05",X"01",X"00",X"02",X"01",X"01",X"05",X"01",X"02",X"1A",X"FF",X"50",X"AA",X"AA",
		X"01",X"FF",X"26",X"01",X"00",X"04",X"01",X"01",X"26",X"FF",X"60",X"AA",X"AA",X"02",X"FF",X"0F",
		X"01",X"FF",X"01",X"01",X"00",X"02",X"01",X"01",X"01",X"02",X"01",X"1F",X"FF",X"30",X"AA",X"AA",
		X"01",X"FE",X"1D",X"01",X"FF",X"02",X"01",X"00",X"02",X"01",X"01",X"02",X"01",X"02",X"0D",X"FF",
		X"28",X"AA",X"AA",X"01",X"FE",X"10",X"01",X"FF",X"03",X"01",X"00",X"02",X"01",X"01",X"03",X"01",
		X"02",X"07",X"01",X"03",X"09",X"00",X"03",X"01",X"00",X"04",X"01",X"FF",X"50",X"AA",X"AA",X"01",
		X"FF",X"26",X"01",X"00",X"04",X"01",X"01",X"26",X"FF",X"30",X"AA",X"AA",X"01",X"FE",X"12",X"01",
		X"FF",X"05",X"01",X"00",X"02",X"01",X"01",X"05",X"01",X"02",X"12",X"FF",X"28",X"AA",X"AA",X"01",
		X"FE",X"10",X"01",X"FF",X"03",X"01",X"00",X"02",X"01",X"01",X"03",X"01",X"02",X"07",X"01",X"03",
		X"09",X"00",X"03",X"01",X"00",X"04",X"01",X"FF",X"38",X"AA",X"AA",X"01",X"FE",X"12",X"01",X"FF",
		X"05",X"01",X"00",X"02",X"01",X"01",X"05",X"01",X"02",X"0A",X"FF",X"50",X"AA",X"AA",X"01",X"FF",
		X"26",X"01",X"00",X"04",X"01",X"01",X"26",X"FF",X"28",X"AA",X"AA",X"01",X"FE",X"13",X"01",X"FF",
		X"04",X"01",X"00",X"02",X"01",X"01",X"04",X"01",X"02",X"0B",X"FF",X"50",X"AA",X"AA",X"01",X"FE",
		X"25",X"01",X"FF",X"02",X"01",X"00",X"02",X"01",X"01",X"02",X"01",X"02",X"25",X"FF",X"30",X"AA",
		X"AA",X"01",X"FE",X"1B",X"01",X"FF",X"04",X"01",X"00",X"02",X"01",X"01",X"04",X"01",X"02",X"0B",
		X"FF",X"50",X"AA",X"AA",X"01",X"FF",X"37",X"01",X"00",X"02",X"01",X"01",X"17",X"FF",X"50",X"AA",
		X"AA",X"01",X"FF",X"26",X"01",X"00",X"04",X"01",X"01",X"26",X"FF",X"B3",X"09",X"C7",X"09",X"D5",
		X"09",X"E9",X"09",X"C8",X"30",X"AA",X"AA",X"01",X"FE",X"1B",X"01",X"FF",X"04",X"01",X"00",X"02",
		X"01",X"01",X"04",X"01",X"02",X"0B",X"FF",X"C8",X"50",X"AA",X"AA",X"01",X"FF",X"37",X"01",X"00",
		X"02",X"01",X"01",X"17",X"FF",X"D0",X"28",X"AA",X"AA",X"01",X"FE",X"13",X"01",X"FF",X"04",X"01",
		X"00",X"02",X"01",X"01",X"04",X"01",X"02",X"0B",X"FF",X"E8",X"40",X"AA",X"AA",X"02",X"FF",X"18",
		X"02",X"01",X"08",X"FF",X"00",X"08",X"02",X"00",X"10",X"01",X"00",X"08",X"01",X"00",X"10",X"01",
		X"00",X"08",X"04",X"00",X"08",X"04",X"00",X"08",X"01",X"00",X"08",X"01",X"00",X"08",X"04",X"00",
		X"08",X"04",X"00",X"08",X"01",X"08",X"02",X"00",X"20",X"02",X"00",X"08",X"01",X"00",X"08",X"01",
		X"00",X"10",X"04",X"08",X"01",X"00",X"10",X"01",X"08",X"04",X"1C",X"01",X"00",X"08",X"02",X"18",
		X"01",X"18",X"02",X"00",X"08",X"02",X"08",X"08",X"00",X"08",X"08",X"00",X"08",X"08",X"00",X"10",
		X"08",X"00",X"10",X"04",X"18",X"01",X"00",X"20",X"04",X"08",X"01",X"FF",X"02",X"57",X"0A",X"67",
		X"0A",X"7B",X"0A",X"99",X"0A",X"AF",X"0A",X"50",X"04",X"20",X"08",X"30",X"04",X"30",X"08",X"10",
		X"01",X"10",X"02",X"30",X"01",X"FF",X"08",X"30",X"02",X"40",X"01",X"30",X"02",X"30",X"01",X"20",
		X"08",X"30",X"01",X"10",X"02",X"20",X"01",X"40",X"04",X"FF",X"02",X"60",X"01",X"10",X"08",X"50",
		X"01",X"40",X"08",X"10",X"04",X"20",X"02",X"20",X"04",X"10",X"02",X"20",X"04",X"10",X"08",X"20",
		X"04",X"20",X"08",X"10",X"04",X"30",X"01",X"FF",X"08",X"20",X"02",X"10",X"04",X"20",X"02",X"10",
		X"04",X"40",X"02",X"10",X"04",X"10",X"08",X"10",X"04",X"60",X"08",X"30",X"04",X"FF",X"02",X"30",
		X"08",X"30",X"04",X"FF",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"20",X"4E",X"21",X"90",X"4A",X"06",X"04",X"CF",X"FD",X"21",X"90",X"4A",X"DD",X"21",X"63",
		X"48",X"DD",X"36",X"01",X"33",X"DD",X"36",X"02",X"B0",X"DD",X"36",X"03",X"01",X"DD",X"36",X"04",
		X"38",X"21",X"AA",X"AA",X"22",X"91",X"4A",X"FD",X"36",X"03",X"04",X"3E",X"23",X"06",X"02",X"FF",
		X"FD",X"21",X"90",X"4A",X"DD",X"21",X"63",X"48",X"FD",X"7E",X"00",X"B7",X"20",X"3B",X"DD",X"7E",
		X"02",X"FE",X"B0",X"20",X"0B",X"3A",X"44",X"48",X"FE",X"4C",X"38",X"04",X"FE",X"A0",X"38",X"DB",
		X"FE",X"A0",X"20",X"0A",X"DD",X"36",X"01",X"B3",X"FD",X"34",X"00",X"C3",X"2B",X"0B",X"FD",X"7E",
		X"03",X"B7",X"20",X"45",X"FD",X"36",X"03",X"04",X"DD",X"7E",X"01",X"1E",X"34",X"FE",X"33",X"28",
		X"02",X"1E",X"33",X"DD",X"73",X"01",X"C3",X"A9",X"0B",X"DD",X"7E",X"02",X"FE",X"B0",X"20",X"0E",
		X"DD",X"36",X"01",X"33",X"DD",X"36",X"00",X"00",X"FD",X"35",X"00",X"C3",X"2B",X"0B",X"FD",X"7E",
		X"03",X"B7",X"20",X"15",X"FD",X"36",X"03",X"04",X"DD",X"7E",X"01",X"1E",X"B4",X"FE",X"B3",X"28",
		X"02",X"1E",X"B3",X"DD",X"73",X"01",X"C3",X"A9",X"0B",X"FD",X"35",X"03",X"2A",X"91",X"4A",X"29",
		X"38",X"06",X"22",X"91",X"4A",X"C3",X"2B",X"0B",X"11",X"00",X"00",X"ED",X"5A",X"22",X"91",X"4A",
		X"01",X"01",X"00",X"FD",X"CB",X"00",X"46",X"20",X"03",X"01",X"FF",X"00",X"DD",X"66",X"02",X"DD",
		X"6E",X"04",X"CD",X"A5",X"91",X"DD",X"74",X"02",X"DD",X"75",X"04",X"DD",X"36",X"00",X"00",X"C3",
		X"2B",X"0B",X"DD",X"36",X"01",X"33",X"DD",X"36",X"00",X"00",X"3E",X"60",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"60",X"4E",X"3E",X"90",X"32",X"98",X"4A",X"21",X"68",X"48",X"22",X"99",X"4A",X"3E",X"23",
		X"06",X"01",X"FF",X"2A",X"D8",X"49",X"7D",X"B4",X"CA",X"73",X"0C",X"2B",X"22",X"D8",X"49",X"3A",
		X"98",X"4A",X"B7",X"28",X"E9",X"06",X"08",X"C5",X"2A",X"99",X"4A",X"7E",X"CB",X"7F",X"20",X"2C",
		X"CB",X"5F",X"20",X"28",X"FE",X"20",X"30",X"24",X"F5",X"11",X"68",X"48",X"B7",X"ED",X"52",X"7D",
		X"CD",X"EA",X"91",X"CD",X"1E",X"92",X"CD",X"83",X"26",X"30",X"03",X"F1",X"18",X"0E",X"F1",X"E5",
		X"E6",X"07",X"CD",X"76",X"95",X"E1",X"01",X"02",X"02",X"CD",X"5C",X"90",X"C1",X"2A",X"99",X"4A",
		X"23",X"22",X"99",X"4A",X"3A",X"98",X"4A",X"3D",X"32",X"98",X"4A",X"CA",X"0E",X"0C",X"10",X"B7",
		X"C3",X"0E",X"0C",X"21",X"01",X"48",X"CB",X"56",X"CB",X"96",X"3E",X"90",X"32",X"98",X"4A",X"21",
		X"68",X"48",X"22",X"99",X"4A",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"98",X"4A",X"B7",X"CA",X"D3",
		X"0C",X"06",X"08",X"C5",X"2A",X"99",X"4A",X"3E",X"88",X"A6",X"20",X"20",X"7E",X"FE",X"20",X"30",
		X"1B",X"11",X"68",X"48",X"B7",X"ED",X"52",X"7D",X"CD",X"EA",X"91",X"CD",X"1E",X"92",X"CD",X"83",
		X"26",X"38",X"09",X"AF",X"1E",X"16",X"01",X"02",X"02",X"CD",X"0C",X"90",X"C1",X"2A",X"99",X"4A",
		X"23",X"22",X"99",X"4A",X"3A",X"98",X"4A",X"3D",X"32",X"98",X"4A",X"CA",X"D3",X"0C",X"10",X"C3",
		X"C3",X"85",X"0C",X"3E",X"60",X"FF",X"21",X"01",X"48",X"CB",X"56",X"CB",X"D6",X"21",X"FB",X"0C",
		X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"CD",X"1D",X"94",X"ED",X"53",X"D8",
		X"49",X"3E",X"13",X"FF",X"3E",X"03",X"01",X"00",X"0C",X"FF",X"C9",X"F0",X"00",X"B4",X"00",X"80",
		X"00",X"B4",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"80",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"A0",X"4E",X"CD",X"3E",X"0E",X"3A",X"A6",X"49",X"CB",X"6F",X"28",X"02",X"1E",X"78",X"16",
		X"3C",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"01",X"48",X"E6",X"03",X"20",X"F4",X"CD",X"42",X"0D",
		X"18",X"EF",X"15",X"20",X"09",X"16",X"3C",X"2A",X"94",X"49",X"23",X"22",X"94",X"49",X"1D",X"C0",
		X"3A",X"A6",X"49",X"CB",X"6F",X"C2",X"D0",X"0D",X"CD",X"3E",X"0E",X"D5",X"21",X"C3",X"0D",X"11",
		X"93",X"49",X"06",X"06",X"CD",X"EF",X"8F",X"1E",X"02",X"3A",X"A6",X"49",X"CB",X"67",X"20",X"28",
		X"21",X"CA",X"0D",X"11",X"8E",X"49",X"06",X"06",X"CD",X"80",X"90",X"1E",X"05",X"FE",X"01",X"20",
		X"17",X"21",X"A6",X"49",X"CB",X"66",X"CB",X"E6",X"2A",X"39",X"48",X"11",X"83",X"A0",X"B7",X"ED",
		X"52",X"28",X"05",X"3E",X"1C",X"CD",X"40",X"03",X"21",X"FC",X"42",X"DD",X"21",X"8E",X"49",X"06",
		X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",X"C4",X"0D",X"11",X"8E",X"49",X"06",X"06",X"CD",X"80",
		X"90",X"D1",X"FE",X"00",X"C0",X"3A",X"A6",X"49",X"CB",X"EF",X"32",X"A6",X"49",X"C9",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"1E",X"78",X"D5",X"21",X"73",X"48",X"16",X"00",X"3A",X"96",X"49",X"5F",X"B7",X"ED",X"52",X"E5",
		X"06",X"0C",X"11",X"0C",X"00",X"CB",X"5E",X"20",X"31",X"19",X"10",X"F9",X"E1",X"E5",X"06",X"0C",
		X"CB",X"DE",X"19",X"10",X"FB",X"E1",X"B7",X"11",X"68",X"48",X"ED",X"52",X"7D",X"CD",X"EA",X"91",
		X"CD",X"1E",X"92",X"06",X"01",X"CD",X"1F",X"0E",X"3A",X"36",X"48",X"CB",X"7F",X"20",X"05",X"3E",
		X"09",X"CD",X"40",X"03",X"21",X"96",X"49",X"34",X"D1",X"C9",X"E1",X"D1",X"1E",X"01",X"C9",X"E5",
		X"C5",X"06",X"0C",X"E5",X"C5",X"01",X"02",X"02",X"3E",X"88",X"1E",X"03",X"CD",X"5C",X"90",X"C1",
		X"E1",X"11",X"40",X"00",X"19",X"10",X"EC",X"C1",X"E1",X"2B",X"2B",X"10",X"E2",X"C9",X"D5",X"3A",
		X"AA",X"49",X"FE",X"05",X"38",X"02",X"3E",X"05",X"3D",X"21",X"53",X"0E",X"16",X"00",X"5F",X"19",
		X"D1",X"5E",X"C9",X"09",X"08",X"08",X"08",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"E0",X"4D",X"3A",X"AB",X"49",X"21",X"0F",X"0F",X"CD",X"10",X"94",X"11",X"8E",X"49",X"01",
		X"06",X"00",X"ED",X"B0",X"CD",X"FC",X"0E",X"3E",X"23",X"06",X"01",X"FF",X"15",X"20",X"F8",X"21",
		X"BE",X"0E",X"3A",X"AB",X"49",X"CD",X"1D",X"94",X"EB",X"11",X"93",X"49",X"06",X"06",X"CD",X"EF",
		X"8F",X"21",X"FC",X"42",X"DD",X"21",X"8E",X"49",X"1E",X"05",X"06",X"06",X"0E",X"00",X"CD",X"1E",
		X"90",X"21",X"F6",X"0E",X"11",X"8E",X"49",X"06",X"06",X"CD",X"80",X"90",X"FE",X"00",X"28",X"02",
		X"18",X"C2",X"3E",X"11",X"FF",X"3E",X"01",X"01",X"0F",X"1D",X"FF",X"3E",X"60",X"FF",X"D1",X"0E",
		X"D7",X"0E",X"DD",X"0E",X"E3",X"0E",X"E9",X"0E",X"EF",X"0E",X"F5",X"0E",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"AB",X"49",X"21",
		X"08",X"0F",X"16",X"00",X"5F",X"19",X"56",X"C9",X"03",X"03",X"03",X"03",X"03",X"02",X"03",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"5E",X"0F",X"D7",X"0F",X"38",X"10",X"B1",X"10",X"1E",X"11",X"9D",X"11",X"4C",X"12",X"14",X"40",
		X"04",X"02",X"09",X"C6",X"40",X"40",X"04",X"02",X"09",X"C6",X"42",X"40",X"04",X"02",X"04",X"04",
		X"41",X"40",X"04",X"02",X"04",X"84",X"42",X"40",X"04",X"0E",X"02",X"0D",X"41",X"40",X"04",X"0A",
		X"02",X"44",X"41",X"40",X"03",X"02",X"0C",X"4A",X"41",X"40",X"03",X"02",X"0C",X"4A",X"42",X"40",
		X"03",X"06",X"02",X"8A",X"41",X"40",X"03",X"06",X"02",X"94",X"41",X"40",X"00",X"02",X"03",X"C1",
		X"41",X"40",X"00",X"02",X"02",X"D6",X"41",X"40",X"00",X"02",X"04",X"C6",X"41",X"40",X"00",X"02",
		X"01",X"CC",X"41",X"40",X"00",X"02",X"02",X"CF",X"41",X"40",X"04",X"02",X"02",X"4D",X"42",X"80",
		X"04",X"01",X"01",X"A7",X"41",X"81",X"04",X"01",X"01",X"8B",X"42",X"82",X"04",X"01",X"01",X"2B",
		X"41",X"83",X"04",X"01",X"01",X"16",X"42",X"10",X"40",X"00",X"02",X"02",X"D6",X"41",X"40",X"00",
		X"02",X"02",X"CB",X"41",X"40",X"00",X"02",X"03",X"C1",X"41",X"40",X"14",X"0E",X"02",X"04",X"41",
		X"40",X"14",X"02",X"09",X"06",X"41",X"40",X"14",X"0E",X"02",X"0D",X"41",X"40",X"14",X"02",X"07",
		X"86",X"42",X"40",X"05",X"02",X"02",X"4B",X"41",X"40",X"05",X"0A",X"02",X"49",X"41",X"40",X"05",
		X"02",X"0B",X"4B",X"42",X"40",X"05",X"0A",X"02",X"54",X"41",X"40",X"05",X"02",X"05",X"4F",X"41",
		X"80",X"04",X"01",X"01",X"0C",X"42",X"81",X"04",X"01",X"01",X"CE",X"42",X"82",X"04",X"01",X"01",
		X"EE",X"40",X"83",X"04",X"01",X"01",X"B6",X"41",X"14",X"40",X"00",X"02",X"02",X"D6",X"41",X"40",
		X"00",X"02",X"02",X"C8",X"41",X"40",X"00",X"02",X"03",X"C1",X"41",X"40",X"03",X"06",X"06",X"90",
		X"41",X"40",X"04",X"06",X"02",X"D2",X"41",X"40",X"04",X"02",X"0A",X"4A",X"41",X"40",X"14",X"02",
		X"07",X"06",X"42",X"40",X"14",X"0A",X"02",X"C6",X"40",X"40",X"14",X"02",X"07",X"C8",X"40",X"40",
		X"14",X"08",X"02",X"0D",X"41",X"40",X"04",X"02",X"0A",X"4A",X"42",X"40",X"05",X"02",X"09",X"84",
		X"41",X"40",X"05",X"0A",X"02",X"C4",X"41",X"40",X"05",X"02",X"09",X"C6",X"42",X"40",X"05",X"06",
		X"02",X"0D",X"42",X"40",X"04",X"08",X"02",X"8A",X"41",X"80",X"04",X"01",X"01",X"65",X"41",X"81",
		X"04",X"01",X"01",X"8B",X"42",X"82",X"04",X"01",X"01",X"AA",X"40",X"83",X"04",X"01",X"01",X"16",
		X"42",X"12",X"40",X"03",X"06",X"06",X"D0",X"41",X"40",X"04",X"06",X"06",X"4E",X"41",X"40",X"03",
		X"02",X"02",X"D0",X"41",X"40",X"02",X"06",X"06",X"C8",X"40",X"40",X"05",X"06",X"06",X"C8",X"41",
		X"40",X"03",X"0A",X"06",X"44",X"41",X"40",X"05",X"03",X"02",X"C8",X"41",X"40",X"00",X"02",X"02",
		X"12",X"42",X"40",X"00",X"02",X"02",X"90",X"41",X"40",X"00",X"02",X"02",X"0A",X"41",X"40",X"00",
		X"02",X"02",X"0A",X"42",X"40",X"00",X"06",X"02",X"86",X"41",X"40",X"00",X"02",X"02",X"D6",X"41",
		X"40",X"00",X"02",X"03",X"C1",X"41",X"80",X"04",X"01",X"01",X"25",X"41",X"81",X"04",X"01",X"01",
		X"8D",X"42",X"82",X"04",X"01",X"01",X"AD",X"40",X"83",X"04",X"01",X"01",X"B5",X"41",X"15",X"40",
		X"03",X"10",X"02",X"94",X"40",X"40",X"03",X"10",X"02",X"91",X"40",X"40",X"03",X"10",X"02",X"8E",
		X"40",X"40",X"03",X"16",X"02",X"8A",X"40",X"40",X"03",X"18",X"02",X"87",X"40",X"40",X"03",X"14",
		X"02",X"04",X"41",X"40",X"00",X"02",X"02",X"D6",X"41",X"40",X"00",X"02",X"01",X"53",X"41",X"40",
		X"00",X"02",X"01",X"53",X"42",X"40",X"00",X"02",X"01",X"D0",X"40",X"40",X"00",X"02",X"01",X"D0",
		X"41",X"40",X"00",X"02",X"02",X"4C",X"41",X"40",X"00",X"02",X"01",X"C9",X"41",X"40",X"00",X"02",
		X"01",X"C9",X"42",X"40",X"00",X"02",X"01",X"46",X"41",X"40",X"00",X"02",X"01",X"46",X"42",X"40",
		X"00",X"02",X"03",X"C1",X"41",X"80",X"04",X"01",X"01",X"86",X"42",X"81",X"04",X"01",X"01",X"2C",
		X"41",X"82",X"04",X"01",X"01",X"6F",X"40",X"83",X"04",X"01",X"01",X"16",X"42",X"1D",X"FF",X"0E",
		X"14",X"02",X"03",X"41",X"FF",X"0E",X"10",X"02",X"46",X"41",X"FF",X"0E",X"0E",X"02",X"09",X"41",
		X"FF",X"0E",X"0E",X"02",X"CC",X"40",X"FF",X"0E",X"0E",X"02",X"8F",X"40",X"FF",X"0E",X"0C",X"02",
		X"12",X"41",X"FE",X"0E",X"02",X"01",X"04",X"41",X"FE",X"0E",X"02",X"01",X"44",X"43",X"FE",X"0E",
		X"02",X"01",X"47",X"41",X"FE",X"0E",X"02",X"01",X"07",X"43",X"FE",X"0E",X"02",X"01",X"0A",X"41",
		X"FE",X"0E",X"02",X"01",X"8A",X"42",X"FE",X"0E",X"02",X"01",X"CD",X"40",X"FE",X"0E",X"02",X"01",
		X"4D",X"42",X"FE",X"0E",X"02",X"01",X"90",X"40",X"FE",X"0E",X"02",X"01",X"10",X"42",X"FE",X"0E",
		X"02",X"01",X"13",X"41",X"FE",X"0E",X"02",X"01",X"53",X"42",X"1F",X"00",X"02",X"17",X"C1",X"41",
		X"FE",X"1E",X"02",X"02",X"C3",X"41",X"FE",X"1E",X"02",X"02",X"C6",X"41",X"FE",X"1E",X"02",X"02",
		X"C9",X"41",X"FE",X"1E",X"02",X"02",X"CC",X"41",X"FE",X"1E",X"02",X"02",X"CF",X"41",X"FE",X"1E",
		X"02",X"02",X"D2",X"41",X"80",X"04",X"01",X"01",X"05",X"42",X"81",X"04",X"01",X"01",X"0B",X"42",
		X"82",X"04",X"01",X"01",X"B1",X"41",X"83",X"04",X"01",X"01",X"15",X"42",X"1F",X"FF",X"0E",X"05",
		X"01",X"81",X"42",X"FF",X"0E",X"0C",X"01",X"E2",X"41",X"FF",X"0E",X"10",X"01",X"A3",X"41",X"FF",
		X"0E",X"0F",X"01",X"C4",X"41",X"FF",X"0E",X"0F",X"01",X"E5",X"41",X"FF",X"0E",X"10",X"01",X"C6",
		X"41",X"FF",X"0E",X"15",X"01",X"27",X"41",X"FF",X"0E",X"14",X"01",X"28",X"41",X"FF",X"0E",X"15",
		X"01",X"09",X"41",X"FF",X"0E",X"15",X"01",X"EA",X"40",X"FF",X"0E",X"15",X"01",X"CB",X"40",X"FF",
		X"0E",X"15",X"01",X"AC",X"40",X"FF",X"0E",X"14",X"01",X"6D",X"40",X"FF",X"0E",X"12",X"01",X"6E",
		X"40",X"FF",X"0E",X"0F",X"01",X"4F",X"40",X"FF",X"0E",X"0E",X"01",X"50",X"40",X"FF",X"0E",X"0D",
		X"01",X"71",X"40",X"FF",X"0E",X"0C",X"01",X"92",X"40",X"FF",X"0E",X"0D",X"01",X"B3",X"40",X"FF",
		X"0E",X"0C",X"01",X"D4",X"40",X"FF",X"0E",X"09",X"01",X"55",X"41",X"FF",X"0E",X"09",X"01",X"76",
		X"41",X"FE",X"0E",X"02",X"04",X"D4",X"41",X"FE",X"0E",X"02",X"06",X"0E",X"41",X"FE",X"0E",X"02",
		X"06",X"08",X"42",X"FE",X"0E",X"02",X"04",X"C4",X"42",X"FE",X"0E",X"02",X"03",X"C1",X"41",X"80",
		X"04",X"01",X"01",X"06",X"43",X"81",X"04",X"01",X"01",X"EB",X"41",X"82",X"04",X"01",X"01",X"F2",
		X"40",X"83",X"04",X"01",X"01",X"B6",X"41",X"1C",X"99",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",
		X"1C",X"04",X"FD",X"1E",X"D2",X"18",X"F3",X"1F",X"1D",X"1C",X"95",X"03",X"FB",X"1F",X"00",X"00",
		X"F9",X"1F",X"1C",X"05",X"1F",X"1E",X"F7",X"1F",X"F4",X"1F",X"F2",X"1E",X"1D",X"1C",X"94",X"03",
		X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"05",X"1F",X"1E",X"F8",X"1F",X"F5",X"1F",X"F2",X"1E",
		X"1E",X"1C",X"94",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"05",X"1F",X"1E",X"D3",X"18",
		X"F6",X"1F",X"F1",X"1E",X"F0",X"1E",X"94",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"02",
		X"1F",X"1E",X"1F",X"1E",X"97",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"02",X"1F",X"1E",
		X"1E",X"1E",X"97",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"98",X"03",
		X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"98",X"03",X"FB",X"1F",X"00",X"00",
		X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"98",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"01",
		X"1F",X"1E",X"98",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"98",X"03",
		X"FC",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"97",X"04",X"1F",X"1E",X"00",X"00",
		X"00",X"00",X"F9",X"1F",X"1C",X"01",X"1F",X"1E",X"97",X"04",X"1F",X"1E",X"00",X"00",X"00",X"00",
		X"F9",X"1F",X"1C",X"98",X"04",X"1F",X"1E",X"00",X"00",X"00",X"00",X"F9",X"1F",X"1C",X"98",X"04",
		X"1F",X"1E",X"00",X"00",X"00",X"00",X"F9",X"1F",X"1C",X"98",X"04",X"1F",X"1E",X"00",X"00",X"00",
		X"00",X"F9",X"1F",X"1C",X"98",X"04",X"1F",X"1E",X"00",X"00",X"00",X"00",X"F9",X"1F",X"1C",X"97",
		X"05",X"FD",X"1E",X"1F",X"1E",X"00",X"00",X"00",X"00",X"F9",X"1F",X"1C",X"90",X"0C",X"FD",X"1E",
		X"1F",X"1E",X"1F",X"1E",X"1F",X"1E",X"1F",X"1E",X"1F",X"1E",X"1F",X"1E",X"1F",X"1E",X"1E",X"1E",
		X"FA",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"90",X"02",X"1F",X"1E",X"1E",X"1E",X"87",X"03",X"FB",
		X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"90",X"0C",X"1F",X"1E",X"00",X"00",X"5F",X"19",X"3E",X"1B",
		X"5F",X"1B",X"2E",X"1C",X"1D",X"1B",X"00",X"00",X"00",X"00",X"FB",X"1F",X"00",X"00",X"F9",X"1F",
		X"1C",X"90",X"0C",X"1F",X"1E",X"00",X"00",X"5E",X"19",X"3F",X"1B",X"5E",X"1B",X"3D",X"1C",X"1E",
		X"1B",X"00",X"00",X"00",X"00",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"90",X"0C",X"1F",X"1E",
		X"00",X"00",X"5F",X"19",X"5F",X"1B",X"3E",X"1B",X"2E",X"1C",X"2E",X"1C",X"1D",X"1B",X"00",X"00",
		X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"90",X"0C",X"1F",X"1E",X"5F",X"1D",X"D2",X"1A",X"D0",
		X"1D",X"3F",X"1B",X"2F",X"1C",X"2F",X"1C",X"1F",X"1B",X"1D",X"1B",X"FB",X"1F",X"00",X"00",X"F9",
		X"1F",X"1C",X"90",X"0C",X"5E",X"1D",X"5E",X"1D",X"D3",X"1A",X"D1",X"1D",X"3E",X"1B",X"2F",X"1C",
		X"2F",X"1C",X"1F",X"1B",X"1E",X"1B",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"1C",X"92",X"0A",X"5E",
		X"19",X"5E",X"1B",X"3F",X"1B",X"3D",X"1C",X"3D",X"1C",X"1E",X"1B",X"00",X"00",X"FB",X"1F",X"00",
		X"00",X"F9",X"1F",X"1C",X"99",X"03",X"FB",X"1F",X"00",X"00",X"F9",X"1F",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"3A",X"A4",X"49",X"B7",X"20",X"45",X"3A",X"80",X"50",X"2F",X"E6",X"0C",X"28",X"31",X"CB",X"3F",
		X"CB",X"3F",X"3D",X"21",X"22",X"91",X"CD",X"1D",X"94",X"EB",X"3A",X"A6",X"49",X"FE",X"04",X"30",
		X"1E",X"CD",X"10",X"94",X"E5",X"DD",X"E1",X"21",X"38",X"41",X"1E",X"17",X"06",X"06",X"0E",X"00",
		X"CD",X"1E",X"90",X"DD",X"21",X"FE",X"15",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"10",X"FF",X"DD",
		X"21",X"C2",X"15",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"10",X"FF",X"21",X"00",X"4B",X"06",X"06",
		X"CF",X"3E",X"01",X"32",X"01",X"4B",X"11",X"05",X"4B",X"21",X"8D",X"49",X"06",X"06",X"CD",X"EF",
		X"8F",X"0E",X"00",X"06",X"05",X"11",X"01",X"4B",X"DD",X"21",X"89",X"40",X"D5",X"DD",X"E5",X"1A",
		X"B9",X"28",X"40",X"C5",X"F5",X"3E",X"1B",X"CD",X"40",X"03",X"F1",X"C1",X"0E",X"FF",X"C5",X"21",
		X"1B",X"16",X"CD",X"1D",X"94",X"EB",X"01",X"03",X"07",X"C5",X"DD",X"E5",X"7E",X"23",X"DD",X"77",
		X"00",X"DD",X"E5",X"11",X"00",X"04",X"DD",X"19",X"DD",X"36",X"00",X"05",X"DD",X"E1",X"DD",X"23",
		X"10",X"EA",X"3E",X"23",X"06",X"03",X"FF",X"DD",X"E1",X"11",X"20",X"00",X"DD",X"19",X"C1",X"0D",
		X"20",X"D7",X"C1",X"DD",X"E1",X"11",X"A0",X"00",X"DD",X"19",X"D1",X"13",X"05",X"C2",X"5C",X"15",
		X"3A",X"A4",X"49",X"B7",X"DD",X"21",X"E2",X"15",X"28",X"04",X"DD",X"21",X"EF",X"15",X"CD",X"0A",
		X"8F",X"C9",X"00",X"0D",X"55",X"41",X"00",X"04",X"59",X"4F",X"55",X"52",X"20",X"50",X"52",X"45",
		X"53",X"53",X"49",X"4E",X"47",X"07",X"B3",X"41",X"00",X"04",X"47",X"4F",X"41",X"4C",X"20",X"49",
		X"53",X"00",X"00",X"06",X"E6",X"42",X"00",X"04",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"00",
		X"08",X"66",X"42",X"00",X"04",X"54",X"4F",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",X"00",X"0B",
		X"5A",X"41",X"00",X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4C",X"49",X"56",X"45",X"53",X"06",
		X"18",X"42",X"00",X"00",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"2F",X"16",X"44",X"16",X"59",
		X"16",X"6E",X"16",X"83",X"16",X"98",X"16",X"AD",X"16",X"C2",X"16",X"D7",X"16",X"EC",X"16",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"1F",
		X"1F",X"00",X"1F",X"00",X"00",X"00",X"1F",X"1F",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",
		X"00",X"1F",X"00",X"00",X"1F",X"1F",X"00",X"00",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",
		X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"00",X"00",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",
		X"00",X"1F",X"00",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",
		X"00",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"1F",
		X"1F",X"1F",X"1F",X"1F",X"00",X"00",X"1F",X"00",X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",
		X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"11",X"0E",X"48",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"03",X"11",X"14",X"48",X"06",X"1E",X"21",
		X"00",X"4C",X"0E",X"01",X"C5",X"E5",X"D5",X"06",X"06",X"CD",X"80",X"90",X"D1",X"E1",X"C1",X"FE",
		X"02",X"28",X"0A",X"C5",X"01",X"08",X"00",X"09",X"C1",X"0C",X"10",X"E8",X"C9",X"79",X"F5",X"FE",
		X"1E",X"28",X"19",X"3E",X"1E",X"91",X"21",X"08",X"00",X"3D",X"28",X"06",X"01",X"08",X"00",X"09",
		X"18",X"F7",X"E5",X"C1",X"21",X"E7",X"4C",X"11",X"EF",X"4C",X"ED",X"B8",X"F1",X"F5",X"3D",X"21",
		X"00",X"4C",X"4F",X"87",X"87",X"87",X"06",X"00",X"4F",X"09",X"11",X"0E",X"48",X"3A",X"01",X"48",
		X"CB",X"6F",X"28",X"03",X"11",X"14",X"48",X"EB",X"01",X"06",X"00",X"ED",X"B0",X"EB",X"3A",X"A8",
		X"49",X"77",X"23",X"3A",X"A9",X"49",X"77",X"DD",X"21",X"5E",X"18",X"CD",X"0A",X"8F",X"DD",X"21",
		X"7D",X"18",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"30",X"FF",X"F1",X"F5",X"21",X"00",X"01",X"22",
		X"00",X"4B",X"21",X"00",X"4C",X"FE",X"0B",X"38",X"14",X"11",X"50",X"00",X"19",X"D6",X"0A",X"E5",
		X"2A",X"00",X"4B",X"11",X"01",X"00",X"19",X"22",X"00",X"4B",X"E1",X"18",X"E8",X"CD",X"FA",X"17",
		X"F1",X"FE",X"0B",X"38",X"04",X"D6",X"0A",X"18",X"F8",X"21",X"D6",X"44",X"3D",X"28",X"04",X"2B",
		X"2B",X"18",X"F9",X"06",X"0A",X"C5",X"E5",X"06",X"13",X"36",X"05",X"CD",X"79",X"90",X"10",X"F9",
		X"3E",X"23",X"06",X"10",X"FF",X"E1",X"E5",X"06",X"13",X"36",X"02",X"CD",X"79",X"90",X"10",X"F9",
		X"3E",X"23",X"06",X"08",X"FF",X"E1",X"C1",X"10",X"DC",X"C9",X"E5",X"DD",X"E1",X"21",X"F6",X"40",
		X"06",X"0A",X"C5",X"DD",X"E5",X"E5",X"DD",X"21",X"00",X"4B",X"1E",X"04",X"06",X"02",X"0E",X"00",
		X"CD",X"1E",X"90",X"E1",X"DD",X"E1",X"DD",X"E5",X"E5",X"01",X"C0",X"00",X"09",X"1E",X"17",X"06",
		X"06",X"0E",X"00",X"CD",X"1E",X"90",X"E1",X"DD",X"E1",X"DD",X"E5",X"E5",X"01",X"00",X"02",X"09",
		X"01",X"06",X"00",X"DD",X"09",X"1E",X"00",X"06",X"02",X"0E",X"00",X"CD",X"1E",X"90",X"3E",X"23",
		X"06",X"02",X"FF",X"11",X"01",X"4B",X"21",X"5D",X"18",X"06",X"02",X"CD",X"DA",X"8F",X"E1",X"DD",
		X"E1",X"2B",X"2B",X"01",X"08",X"00",X"DD",X"09",X"C1",X"10",X"A7",X"C9",X"00",X"01",X"00",X"18",
		X"9C",X"40",X"00",X"05",X"54",X"4F",X"44",X"41",X"59",X"3C",X"53",X"20",X"48",X"49",X"3B",X"53",
		X"43",X"4F",X"52",X"45",X"20",X"42",X"45",X"53",X"54",X"20",X"33",X"30",X"00",X"00",X"05",X"D8",
		X"40",X"00",X"04",X"4F",X"52",X"44",X"45",X"52",X"05",X"D8",X"41",X"00",X"17",X"53",X"43",X"4F",
		X"52",X"45",X"05",X"D8",X"42",X"00",X"00",X"52",X"4F",X"55",X"4E",X"44",X"00",X"FF",X"FF",X"FF",
		X"31",X"60",X"4F",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"0F",X"3E",X"05",X"32",X"AB",X"49",X"AF",
		X"32",X"E0",X"4A",X"21",X"39",X"1F",X"22",X"E2",X"4A",X"3E",X"1E",X"CD",X"40",X"03",X"DD",X"21",
		X"2E",X"1F",X"CD",X"0A",X"8F",X"DD",X"21",X"16",X"1F",X"CD",X"0A",X"8F",X"3A",X"AB",X"49",X"3C",
		X"C6",X"30",X"21",X"52",X"42",X"77",X"CB",X"D4",X"36",X"17",X"3E",X"23",X"06",X"40",X"FF",X"CD",
		X"5B",X"35",X"21",X"50",X"0F",X"3A",X"AB",X"49",X"CD",X"1D",X"94",X"D5",X"FD",X"E1",X"FD",X"46",
		X"00",X"FD",X"23",X"C5",X"FD",X"7E",X"00",X"FD",X"23",X"FD",X"5E",X"00",X"FD",X"23",X"FD",X"4E",
		X"00",X"FD",X"23",X"FD",X"46",X"00",X"FD",X"23",X"FD",X"6E",X"00",X"FD",X"23",X"FD",X"66",X"00",
		X"FD",X"23",X"CD",X"4A",X"90",X"C1",X"10",X"DB",X"21",X"40",X"40",X"FD",X"21",X"07",X"13",X"FD",
		X"7E",X"00",X"FD",X"23",X"B7",X"28",X"37",X"4F",X"FD",X"46",X"00",X"FD",X"23",X"CB",X"78",X"CB",
		X"B8",X"20",X"18",X"FD",X"7E",X"00",X"FD",X"23",X"FD",X"5E",X"00",X"FD",X"23",X"77",X"CB",X"D4",
		X"73",X"CB",X"94",X"23",X"0D",X"28",X"0C",X"10",X"EA",X"18",X"DD",X"23",X"0D",X"28",X"04",X"10",
		X"FA",X"18",X"D5",X"7D",X"E6",X"E0",X"6F",X"11",X"20",X"00",X"19",X"C3",X"1F",X"19",X"3E",X"04",
		X"01",X"00",X"96",X"FF",X"3E",X"02",X"01",X"00",X"0B",X"FF",X"21",X"FE",X"1E",X"11",X"00",X"4B",
		X"01",X"18",X"00",X"ED",X"B0",X"3A",X"AB",X"49",X"21",X"1D",X"1E",X"CD",X"16",X"94",X"11",X"02",
		X"4B",X"01",X"04",X"00",X"ED",X"B0",X"21",X"E0",X"49",X"06",X"20",X"CF",X"FD",X"21",X"E0",X"49",
		X"DD",X"21",X"40",X"48",X"DD",X"36",X"01",X"0E",X"DD",X"36",X"02",X"80",X"DD",X"36",X"03",X"81",
		X"DD",X"36",X"04",X"F8",X"FD",X"36",X"02",X"D6",X"FD",X"36",X"03",X"D6",X"3E",X"17",X"CD",X"40",
		X"03",X"3E",X"03",X"01",X"60",X"0E",X"FF",X"DD",X"36",X"00",X"00",X"3E",X"23",X"06",X"02",X"FF",
		X"CD",X"A1",X"1E",X"3E",X"50",X"DD",X"BE",X"04",X"D2",X"78",X"1B",X"3A",X"1A",X"48",X"E6",X"01",
		X"C4",X"6C",X"1A",X"CD",X"39",X"1E",X"30",X"DF",X"CD",X"66",X"2E",X"CD",X"24",X"94",X"21",X"1C",
		X"1A",X"16",X"00",X"5F",X"19",X"7E",X"47",X"FE",X"02",X"20",X"0B",X"3E",X"F8",X"DD",X"BE",X"04",
		X"78",X"20",X"03",X"3E",X"04",X"47",X"FD",X"BE",X"01",X"CA",X"3C",X"1A",X"DD",X"7E",X"02",X"E6",
		X"07",X"C2",X"3C",X"1A",X"DD",X"7E",X"04",X"E6",X"07",X"C2",X"3C",X"1A",X"78",X"FE",X"04",X"20",
		X"10",X"DD",X"36",X"01",X"0E",X"FD",X"36",X"01",X"04",X"C3",X"B7",X"19",X"00",X"03",X"01",X"02",
		X"04",X"C5",X"CD",X"A5",X"1A",X"C1",X"C2",X"3C",X"1A",X"FD",X"70",X"01",X"78",X"21",X"74",X"1B",
		X"16",X"00",X"5F",X"19",X"7E",X"DD",X"77",X"01",X"FD",X"36",X"04",X"00",X"DD",X"7E",X"02",X"E6",
		X"07",X"C2",X"55",X"1A",X"DD",X"7E",X"04",X"E6",X"07",X"C2",X"55",X"1A",X"FD",X"7E",X"01",X"CD",
		X"A5",X"1A",X"C2",X"5F",X"1A",X"3E",X"04",X"FD",X"BE",X"01",X"28",X"03",X"CD",X"F8",X"2D",X"3E",
		X"04",X"FD",X"BE",X"01",X"28",X"03",X"CD",X"49",X"2E",X"C3",X"B7",X"19",X"DD",X"7E",X"02",X"C6",
		X"F4",X"5F",X"C6",X"18",X"57",X"DD",X"7E",X"04",X"C6",X"F4",X"6F",X"C6",X"18",X"67",X"DD",X"E5",
		X"DD",X"21",X"45",X"48",X"06",X"06",X"DD",X"7E",X"02",X"BB",X"38",X"0D",X"BA",X"30",X"0A",X"DD",
		X"7E",X"04",X"BD",X"38",X"04",X"BC",X"DA",X"A3",X"1C",X"C5",X"01",X"05",X"00",X"DD",X"09",X"C1",
		X"10",X"E4",X"DD",X"E1",X"C9",X"F5",X"47",X"3A",X"AB",X"49",X"FE",X"06",X"20",X"1E",X"CB",X"40",
		X"28",X"1A",X"DD",X"7E",X"04",X"FE",X"E0",X"CA",X"CC",X"1A",X"FE",X"C0",X"CA",X"CC",X"1A",X"FE",
		X"90",X"CA",X"CC",X"1A",X"FE",X"60",X"CA",X"CC",X"1A",X"B7",X"F1",X"C9",X"3A",X"AB",X"49",X"21",
		X"2C",X"1B",X"FE",X"05",X"38",X"0A",X"21",X"44",X"1B",X"FE",X"05",X"28",X"03",X"21",X"5C",X"1B",
		X"F1",X"CD",X"10",X"94",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"E5",X"D5",X"C5",X"DD",
		X"66",X"02",X"DD",X"6E",X"04",X"CD",X"1E",X"92",X"C1",X"D1",X"19",X"3A",X"AB",X"49",X"FE",X"05",
		X"38",X"18",X"3E",X"00",X"E5",X"B6",X"23",X"10",X"FC",X"E1",X"0D",X"28",X"05",X"11",X"20",X"00",
		X"19",X"B6",X"E1",X"47",X"AE",X"C8",X"23",X"78",X"AE",X"C9",X"3E",X"FF",X"E5",X"A6",X"23",X"10",
		X"FC",X"E1",X"0D",X"28",X"ED",X"11",X"20",X"00",X"19",X"A6",X"18",X"E6",X"02",X"01",X"02",X"00",
		X"40",X"40",X"01",X"02",X"40",X"00",X"40",X"40",X"02",X"01",X"FF",X"FF",X"40",X"40",X"01",X"02",
		X"E0",X"FF",X"40",X"40",X"02",X"01",X"00",X"00",X"1F",X"FE",X"01",X"02",X"40",X"00",X"1F",X"FE",
		X"02",X"01",X"FF",X"FF",X"1F",X"FE",X"01",X"02",X"E0",X"FF",X"1F",X"FE",X"02",X"01",X"00",X"00",
		X"FE",X"FE",X"01",X"02",X"40",X"00",X"FE",X"FF",X"02",X"01",X"FF",X"FF",X"FE",X"FE",X"01",X"02",
		X"E0",X"FF",X"FE",X"FF",X"0C",X"08",X"0A",X"88",X"3E",X"13",X"FF",X"3E",X"23",X"06",X"02",X"FF",
		X"CD",X"A1",X"1E",X"3E",X"38",X"DD",X"BE",X"04",X"28",X"0E",X"CD",X"39",X"1E",X"30",X"EC",X"CD",
		X"76",X"1E",X"DD",X"36",X"00",X"00",X"18",X"E3",X"3E",X"23",X"06",X"02",X"FF",X"3E",X"90",X"DD",
		X"BE",X"02",X"28",X"0E",X"CD",X"39",X"1E",X"30",X"EF",X"CD",X"8E",X"1E",X"DD",X"36",X"00",X"00",
		X"18",X"E6",X"DD",X"36",X"01",X"32",X"DD",X"36",X"00",X"00",X"3E",X"23",X"06",X"01",X"FF",X"3A",
		X"65",X"48",X"FE",X"A0",X"20",X"F4",X"3E",X"80",X"CD",X"40",X"03",X"3E",X"12",X"FF",X"3E",X"14",
		X"FF",X"21",X"45",X"48",X"06",X"1E",X"CF",X"11",X"45",X"48",X"21",X"9E",X"1C",X"01",X"05",X"00",
		X"ED",X"B0",X"11",X"E1",X"49",X"21",X"4E",X"1E",X"01",X"28",X"00",X"ED",X"B0",X"3E",X"80",X"32",
		X"E0",X"49",X"3E",X"0A",X"CD",X"40",X"03",X"3E",X"23",X"06",X"02",X"FF",X"3A",X"22",X"48",X"CB",
		X"7F",X"CA",X"53",X"1D",X"FD",X"21",X"E0",X"49",X"FD",X"7E",X"00",X"B7",X"CA",X"53",X"1D",X"FD",
		X"35",X"00",X"FD",X"23",X"06",X"08",X"C5",X"FD",X"7E",X"02",X"B7",X"28",X"3A",X"FD",X"35",X"02",
		X"11",X"05",X"00",X"FD",X"19",X"C1",X"10",X"EE",X"FD",X"7E",X"00",X"CB",X"BF",X"B7",X"20",X"21",
		X"3E",X"00",X"FD",X"CB",X"00",X"7E",X"FD",X"CB",X"00",X"BE",X"20",X"06",X"FD",X"CB",X"00",X"FE",
		X"3E",X"1F",X"32",X"46",X"48",X"AF",X"32",X"45",X"48",X"3E",X"0C",X"FD",X"B6",X"00",X"FD",X"77",
		X"00",X"FD",X"35",X"00",X"C3",X"F7",X"1B",X"FD",X"7E",X"03",X"CB",X"BF",X"FD",X"77",X"02",X"FD",
		X"7E",X"04",X"FD",X"CB",X"03",X"7E",X"28",X"12",X"FE",X"19",X"28",X"12",X"FD",X"CB",X"03",X"FE",
		X"D6",X"04",X"FE",X"1D",X"20",X"14",X"D6",X"04",X"18",X"10",X"FE",X"25",X"28",X"EE",X"FD",X"CB",
		X"03",X"BE",X"C6",X"04",X"FE",X"1D",X"20",X"02",X"C6",X"04",X"FD",X"77",X"04",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"1E",X"0D",X"01",X"02",X"02",X"CD",X"5C",X"90",X"C3",X"20",X"1C",X"00",X"1F",
		X"98",X"10",X"30",X"3E",X"13",X"FF",X"3E",X"14",X"FF",X"21",X"45",X"48",X"06",X"1E",X"CF",X"3E",
		X"80",X"CD",X"40",X"03",X"DD",X"21",X"40",X"48",X"DD",X"36",X"01",X"0F",X"3E",X"13",X"CD",X"40",
		X"03",X"3E",X"23",X"06",X"01",X"FF",X"3E",X"FD",X"DD",X"BE",X"04",X"38",X"0E",X"3E",X"02",X"DD",
		X"86",X"04",X"DD",X"77",X"04",X"DD",X"36",X"00",X"00",X"18",X"E6",X"21",X"8E",X"49",X"06",X"06",
		X"CF",X"3E",X"14",X"CD",X"40",X"03",X"DD",X"36",X"04",X"00",X"DD",X"36",X"01",X"10",X"DD",X"36",
		X"00",X"00",X"3E",X"23",X"06",X"28",X"FF",X"3E",X"14",X"CD",X"40",X"03",X"DD",X"36",X"01",X"17",
		X"DD",X"36",X"00",X"00",X"3E",X"12",X"FF",X"3E",X"40",X"06",X"20",X"FF",X"3E",X"60",X"FF",X"31",
		X"60",X"4F",X"3E",X"14",X"FF",X"3E",X"12",X"FF",X"3E",X"23",X"06",X"05",X"FF",X"3E",X"80",X"CD",
		X"40",X"03",X"DD",X"21",X"40",X"48",X"CD",X"82",X"2A",X"21",X"8E",X"49",X"06",X"06",X"CF",X"AF",
		X"5F",X"01",X"0B",X"03",X"21",X"4E",X"41",X"CD",X"4A",X"90",X"DD",X"21",X"43",X"1D",X"CD",X"0A",
		X"8F",X"18",X"C1",X"00",X"09",X"6F",X"41",X"00",X"17",X"54",X"49",X"4D",X"45",X"20",X"4F",X"56",
		X"45",X"52",X"00",X"21",X"00",X"40",X"01",X"00",X"04",X"7E",X"FE",X"80",X"38",X"07",X"FE",X"84",
		X"30",X"03",X"CD",X"EB",X"1E",X"23",X"0B",X"79",X"B0",X"20",X"EE",X"21",X"4A",X"41",X"AF",X"5F",
		X"01",X"08",X"09",X"CD",X"0C",X"90",X"FD",X"21",X"00",X"4B",X"21",X"71",X"41",X"06",X"04",X"0E",
		X"00",X"C5",X"E5",X"FD",X"7E",X"00",X"B7",X"28",X"67",X"E5",X"79",X"21",X"15",X"1E",X"CD",X"1D",
		X"94",X"7A",X"01",X"01",X"01",X"E1",X"E5",X"CD",X"5C",X"90",X"E1",X"11",X"20",X"00",X"19",X"FD",
		X"36",X"00",X"00",X"FD",X"E5",X"DD",X"E1",X"DD",X"23",X"06",X"05",X"0E",X"00",X"1E",X"00",X"CD",
		X"1E",X"90",X"06",X"06",X"3E",X"0A",X"FD",X"E5",X"FD",X"BE",X"00",X"20",X"04",X"FD",X"36",X"00",
		X"00",X"FD",X"23",X"10",X"F3",X"FD",X"E1",X"FD",X"E5",X"E1",X"11",X"05",X"00",X"19",X"11",X"8D",
		X"49",X"06",X"06",X"CD",X"DA",X"8F",X"21",X"BD",X"41",X"DD",X"21",X"88",X"49",X"1E",X"04",X"06",
		X"06",X"0E",X"00",X"CD",X"1E",X"90",X"3E",X"23",X"06",X"08",X"FF",X"E1",X"2B",X"2B",X"18",X"01",
		X"E1",X"C1",X"0C",X"11",X"06",X"00",X"FD",X"19",X"05",X"C2",X"81",X"1D",X"3A",X"AB",X"49",X"3C",
		X"FE",X"07",X"38",X"01",X"AF",X"32",X"AB",X"49",X"3E",X"23",X"06",X"2D",X"FF",X"3E",X"40",X"06",
		X"10",X"FF",X"3E",X"60",X"FF",X"04",X"83",X"04",X"82",X"04",X"81",X"04",X"80",X"02",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"2A",X"E2",X"49",X"29",X"38",X"04",X"22",
		X"E2",X"49",X"C9",X"F5",X"11",X"00",X"00",X"ED",X"5A",X"22",X"E2",X"49",X"F1",X"C9",X"7A",X"40",
		X"00",X"04",X"19",X"BA",X"40",X"00",X"02",X"19",X"FA",X"40",X"00",X"04",X"19",X"3A",X"41",X"00",
		X"02",X"19",X"7A",X"41",X"00",X"04",X"19",X"BA",X"42",X"00",X"02",X"19",X"FA",X"42",X"00",X"04",
		X"19",X"3A",X"43",X"00",X"02",X"19",X"FD",X"7E",X"01",X"E6",X"07",X"20",X"07",X"CD",X"F8",X"2D",
		X"CD",X"49",X"2E",X"C9",X"DD",X"36",X"01",X"0C",X"FD",X"36",X"01",X"00",X"18",X"EF",X"FD",X"7E",
		X"01",X"E6",X"07",X"FE",X"01",X"28",X"E6",X"DD",X"36",X"01",X"08",X"FD",X"36",X"01",X"01",X"18",
		X"DC",X"DD",X"7E",X"02",X"67",X"E6",X"07",X"C0",X"DD",X"7E",X"04",X"6F",X"E6",X"07",X"C0",X"CD",
		X"1E",X"92",X"11",X"E1",X"FF",X"19",X"0E",X"00",X"7E",X"EB",X"21",X"D1",X"1E",X"06",X"04",X"BE",
		X"23",X"28",X"12",X"10",X"FA",X"0C",X"3E",X"02",X"B9",X"C8",X"EB",X"11",X"60",X"00",X"19",X"18",
		X"E7",X"80",X"81",X"82",X"83",X"21",X"00",X"4B",X"4F",X"D6",X"80",X"2F",X"E6",X"03",X"D5",X"CD",
		X"10",X"94",X"D1",X"36",X"01",X"EB",X"3E",X"0F",X"CD",X"40",X"03",X"3A",X"AB",X"49",X"FE",X"06",
		X"3E",X"00",X"20",X"02",X"3E",X"FF",X"77",X"CB",X"D4",X"36",X"0E",X"CB",X"94",X"C9",X"00",X"0A",
		X"01",X"00",X"00",X"00",X"00",X"0A",X"0A",X"08",X"00",X"00",X"00",X"0A",X"0A",X"06",X"00",X"00",
		X"00",X"0A",X"0A",X"04",X"00",X"00",X"04",X"09",X"97",X"41",X"00",X"00",X"50",X"4C",X"41",X"59",
		X"20",X"47",X"41",X"4D",X"45",X"03",X"D2",X"41",X"00",X"05",X"41",X"43",X"54",X"00",X"00",X"05",
		X"1D",X"43",X"00",X"00",X"20",X"54",X"49",X"4D",X"45",X"00",X"0A",X"00",X"04",X"01",X"06",X"00",
		X"02",X"01",X"0D",X"00",X"0D",X"01",X"05",X"00",X"04",X"01",X"05",X"00",X"03",X"01",X"0D",X"00",
		X"0F",X"08",X"0F",X"00",X"28",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FD",X"21",X"80",X"4A",X"FD",X"CB",X"00",X"7E",
		X"C2",X"93",X"22",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"04",X"CD",X"40",X"03",X"FD",X"CB",X"00",
		X"FE",X"CD",X"A9",X"2E",X"3E",X"16",X"32",X"66",X"48",X"3A",X"E9",X"49",X"E6",X"07",X"FD",X"77",
		X"02",X"FD",X"E5",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"AC",X"91",X"EB",X"21",X"68",X"48",
		X"FD",X"21",X"D0",X"4A",X"06",X"90",X"7E",X"E6",X"70",X"FE",X"10",X"28",X"09",X"23",X"10",X"F6",
		X"FD",X"E1",X"D1",X"C3",X"2A",X"24",X"E5",X"B7",X"ED",X"52",X"E1",X"28",X"04",X"FD",X"23",X"18",
		X"EC",X"CB",X"DE",X"7E",X"E6",X"07",X"21",X"7B",X"26",X"16",X"00",X"3D",X"5F",X"19",X"5E",X"FD",
		X"7E",X"00",X"FD",X"E1",X"FD",X"77",X"03",X"21",X"7F",X"26",X"06",X"00",X"4F",X"09",X"7E",X"DD",
		X"66",X"02",X"DD",X"6E",X"04",X"D5",X"F5",X"CD",X"1E",X"92",X"F1",X"D1",X"01",X"02",X"02",X"CD",
		X"5C",X"90",X"C9",X"FD",X"7E",X"01",X"B7",X"28",X"04",X"FD",X"35",X"01",X"C9",X"FD",X"36",X"01",
		X"01",X"CD",X"C7",X"2E",X"C0",X"C1",X"21",X"01",X"48",X"CB",X"46",X"CB",X"C6",X"3E",X"23",X"06",
		X"05",X"FF",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"1E",X"92",X"01",X"02",X"02",X"1E",X"16",
		X"3E",X"00",X"CD",X"0C",X"90",X"FD",X"7E",X"03",X"F6",X"80",X"FD",X"77",X"00",X"FD",X"7E",X"02",
		X"FD",X"77",X"06",X"FD",X"36",X"03",X"83",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"AC",X"91",
		X"FD",X"75",X"04",X"FD",X"74",X"05",X"CB",X"FE",X"CB",X"9E",X"FD",X"36",X"01",X"00",X"21",X"59",
		X"48",X"06",X"0F",X"CF",X"DD",X"21",X"45",X"48",X"3A",X"42",X"48",X"DD",X"77",X"02",X"3A",X"44",
		X"48",X"DD",X"77",X"04",X"21",X"7B",X"26",X"FD",X"7E",X"06",X"16",X"00",X"3D",X"5F",X"19",X"7E",
		X"DD",X"77",X"03",X"3E",X"02",X"CD",X"93",X"25",X"DD",X"36",X"00",X"01",X"FD",X"36",X"07",X"00",
		X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"81",X"CD",X"40",X"03",X"3E",X"08",X"CD",X"40",X"03",X"AF",
		X"32",X"40",X"48",X"32",X"41",X"48",X"3E",X"23",X"06",X"02",X"FF",X"C3",X"3E",X"23",X"3E",X"23",
		X"06",X"01",X"FF",X"FD",X"21",X"80",X"4A",X"DD",X"21",X"45",X"48",X"CD",X"54",X"23",X"DD",X"36",
		X"00",X"01",X"18",X"EA",X"FD",X"CB",X"03",X"7E",X"28",X"10",X"FD",X"7E",X"03",X"CB",X"BF",X"B7",
		X"20",X"05",X"CD",X"69",X"24",X"18",X"03",X"FD",X"35",X"03",X"FD",X"CB",X"01",X"7E",X"28",X"28",
		X"FD",X"7E",X"02",X"B7",X"28",X"04",X"FD",X"35",X"02",X"C9",X"FD",X"CB",X"01",X"76",X"20",X"0E",
		X"FD",X"CB",X"01",X"F6",X"3E",X"01",X"CD",X"93",X"25",X"FD",X"36",X"02",X"04",X"C9",X"AF",X"FD",
		X"77",X"01",X"3E",X"02",X"CD",X"93",X"25",X"C9",X"CD",X"27",X"26",X"CD",X"5C",X"26",X"CA",X"2A",
		X"24",X"DD",X"7E",X"04",X"FD",X"CB",X"00",X"46",X"28",X"03",X"DD",X"7E",X"02",X"E6",X"0F",X"C0",
		X"DD",X"66",X"02",X"DD",X"6E",X"04",X"3A",X"96",X"49",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",
		X"27",X"C6",X"31",X"BD",X"30",X"59",X"CD",X"AC",X"91",X"FE",X"FF",X"28",X"52",X"CB",X"7F",X"28",
		X"39",X"5F",X"E6",X"70",X"FE",X"40",X"CA",X"1F",X"24",X"FE",X"30",X"7B",X"CA",X"1F",X"24",X"E6",
		X"07",X"B7",X"28",X"3B",X"FD",X"5E",X"06",X"BB",X"28",X"35",X"FD",X"36",X"03",X"88",X"FD",X"75",
		X"04",X"FD",X"74",X"05",X"FD",X"CB",X"01",X"FE",X"FD",X"36",X"07",X"00",X"FD",X"36",X"02",X"04",
		X"AF",X"CD",X"93",X"25",X"3E",X"08",X"CD",X"40",X"03",X"C9",X"CB",X"5F",X"20",X"11",X"5F",X"E6",
		X"70",X"20",X"0C",X"7B",X"57",X"E6",X"07",X"FD",X"5E",X"06",X"BB",X"20",X"02",X"18",X"CB",X"FD",
		X"34",X"07",X"3E",X"03",X"FD",X"BE",X"07",X"C0",X"18",X"CA",X"C1",X"21",X"45",X"48",X"06",X"0A",
		X"CF",X"21",X"80",X"4A",X"06",X"08",X"CF",X"FD",X"21",X"E0",X"49",X"DD",X"21",X"40",X"48",X"FD",
		X"36",X"00",X"00",X"DD",X"36",X"01",X"0E",X"DD",X"36",X"00",X"00",X"3E",X"23",X"06",X"04",X"FF",
		X"21",X"01",X"48",X"CB",X"46",X"CB",X"86",X"21",X"68",X"24",X"CD",X"BA",X"2C",X"C2",X"D5",X"2C",
		X"C3",X"E1",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"FD",X"CB",X"03",X"BE",X"FD",X"6E",X"04",
		X"FD",X"66",X"05",X"7E",X"E6",X"07",X"F5",X"11",X"68",X"48",X"B7",X"ED",X"52",X"7D",X"CD",X"EA",
		X"91",X"CD",X"1E",X"92",X"CD",X"83",X"26",X"30",X"03",X"F1",X"E1",X"C9",X"E5",X"FD",X"7E",X"06",
		X"5F",X"3A",X"01",X"48",X"CB",X"57",X"7B",X"28",X"05",X"CD",X"87",X"95",X"18",X"03",X"CD",X"76",
		X"95",X"E1",X"01",X"02",X"02",X"CD",X"5C",X"90",X"FD",X"7E",X"06",X"3D",X"21",X"2B",X"25",X"CD",
		X"17",X"94",X"5E",X"23",X"56",X"EB",X"F1",X"E5",X"3D",X"5F",X"FD",X"7E",X"06",X"3D",X"F5",X"D5",
		X"D1",X"F1",X"E1",X"93",X"16",X"00",X"B7",X"CA",X"E3",X"24",X"E5",X"F5",X"D5",X"7B",X"D1",X"F1",
		X"CB",X"7F",X"28",X"01",X"15",X"E1",X"87",X"5F",X"87",X"83",X"5F",X"19",X"7A",X"06",X"06",X"CB",
		X"7F",X"28",X"05",X"CD",X"BA",X"2C",X"18",X"24",X"E5",X"11",X"8D",X"49",X"CD",X"EF",X"8F",X"E1",
		X"11",X"13",X"48",X"3A",X"01",X"48",X"CB",X"7F",X"28",X"0C",X"CB",X"6F",X"28",X"03",X"11",X"19",
		X"48",X"06",X"06",X"CD",X"EF",X"8F",X"21",X"68",X"24",X"CD",X"BA",X"2C",X"FD",X"6E",X"04",X"FD",
		X"66",X"05",X"7E",X"E6",X"70",X"FE",X"10",X"20",X"06",X"FD",X"46",X"06",X"B0",X"18",X"05",X"FD",
		X"7E",X"06",X"E6",X"07",X"CB",X"FF",X"77",X"CD",X"90",X"3F",X"C9",X"4A",X"25",X"5C",X"25",X"6E",
		X"25",X"80",X"25",X"00",X"00",X"00",X"04",X"05",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",
		X"02",X"05",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"04",X"05",X"00",X"21",X"DF",X"25",X"B7",X"28",X"0A",X"21",X"F7",X"25",X"FE",X"01",X"28",X"03",
		X"21",X"0F",X"26",X"FD",X"7E",X"00",X"CB",X"BF",X"CD",X"10",X"94",X"4E",X"23",X"46",X"23",X"7E",
		X"23",X"5E",X"23",X"56",X"23",X"E5",X"DD",X"77",X"01",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",
		X"A5",X"91",X"DD",X"74",X"02",X"DD",X"75",X"04",X"D5",X"C1",X"CD",X"A5",X"91",X"DD",X"74",X"07",
		X"DD",X"75",X"09",X"E1",X"7E",X"DD",X"77",X"06",X"DD",X"7E",X"03",X"DD",X"77",X"08",X"C9",X"00",
		X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"A3",
		X"00",X"00",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"00",
		X"F8",X"24",X"00",X"10",X"25",X"08",X"00",X"A6",X"F0",X"00",X"A7",X"00",X"08",X"64",X"00",X"F0",
		X"65",X"F8",X"00",X"26",X"10",X"00",X"27",X"FD",X"7E",X"00",X"CB",X"BF",X"21",X"54",X"26",X"CD",
		X"17",X"94",X"4E",X"23",X"46",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"A5",X"91",X"DD",X"74",
		X"02",X"DD",X"75",X"04",X"DD",X"66",X"07",X"DD",X"6E",X"09",X"CD",X"A5",X"91",X"DD",X"74",X"07",
		X"DD",X"75",X"09",X"C9",X"00",X"FE",X"02",X"00",X"00",X"02",X"FE",X"00",X"FD",X"7E",X"00",X"CB",
		X"BF",X"21",X"73",X"26",X"CD",X"17",X"94",X"7E",X"23",X"DD",X"BE",X"02",X"C8",X"7E",X"DD",X"BE",
		X"04",X"C8",X"C9",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"0E",X"0F",X"10",X"B0",
		X"B8",X"B4",X"BC",X"3A",X"96",X"49",X"B7",X"C8",X"E5",X"CB",X"27",X"67",X"7D",X"E6",X"1F",X"6F",
		X"3E",X"1F",X"95",X"D6",X"06",X"D8",X"BC",X"E1",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"60",X"4F",X"3A",X"01",X"48",X"CB",X"7F",X"28",X"08",X"3A",X"A7",X"49",X"47",X"05",X"CD",
		X"70",X"91",X"CD",X"B6",X"2D",X"21",X"E0",X"49",X"06",X"20",X"CF",X"CD",X"D6",X"2D",X"DD",X"21",
		X"40",X"48",X"DD",X"36",X"01",X"0E",X"DD",X"36",X"02",X"80",X"DD",X"36",X"03",X"81",X"DD",X"36",
		X"04",X"F0",X"3E",X"3C",X"32",X"EC",X"49",X"AF",X"32",X"E0",X"4A",X"21",X"F3",X"09",X"22",X"E2",
		X"4A",X"3E",X"23",X"06",X"02",X"FF",X"FD",X"21",X"E0",X"49",X"DD",X"21",X"40",X"48",X"3A",X"96",
		X"49",X"FE",X"0C",X"CA",X"65",X"2A",X"3A",X"1A",X"48",X"E6",X"01",X"C4",X"F9",X"29",X"3A",X"02",
		X"48",X"CB",X"77",X"28",X"41",X"FD",X"E5",X"FD",X"21",X"A0",X"4A",X"06",X"03",X"FD",X"7E",X"00",
		X"FE",X"02",X"20",X"29",X"FD",X"7E",X"03",X"C6",X"F8",X"57",X"C6",X"50",X"5F",X"DD",X"7E",X"02",
		X"BA",X"38",X"1A",X"BB",X"30",X"17",X"FD",X"7E",X"04",X"C6",X"B8",X"57",X"C6",X"50",X"5F",X"DD",
		X"7E",X"04",X"BA",X"38",X"08",X"BB",X"30",X"05",X"FD",X"E1",X"C3",X"65",X"2A",X"11",X"0A",X"00",
		X"FD",X"19",X"10",X"C9",X"FD",X"E1",X"FD",X"CB",X"00",X"7E",X"CA",X"9B",X"27",X"FD",X"7E",X"00",
		X"CB",X"BF",X"21",X"58",X"27",X"F7",X"18",X"0A",X"79",X"2B",X"08",X"22",X"79",X"2B",X"79",X"2B",
		X"01",X"2B",X"DD",X"21",X"40",X"48",X"FD",X"21",X"E0",X"49",X"FD",X"CB",X"0A",X"76",X"28",X"12",
		X"FD",X"7E",X"0F",X"B7",X"28",X"05",X"FD",X"35",X"0F",X"18",X"07",X"FD",X"CB",X"0A",X"B6",X"CD",
		X"D6",X"2D",X"DD",X"7E",X"01",X"FD",X"77",X"05",X"DD",X"7E",X"02",X"FD",X"77",X"06",X"DD",X"7E",
		X"04",X"FD",X"77",X"07",X"DD",X"36",X"00",X"00",X"C3",X"E1",X"26",X"2A",X"E2",X"49",X"29",X"38",
		X"06",X"22",X"E2",X"49",X"C3",X"62",X"27",X"11",X"00",X"00",X"ED",X"5A",X"22",X"E2",X"49",X"CD",
		X"66",X"2E",X"CD",X"24",X"94",X"21",X"BB",X"27",X"F7",X"18",X"0A",X"52",X"28",X"14",X"29",X"B2",
		X"28",X"76",X"29",X"D6",X"29",X"3E",X"0F",X"DD",X"A6",X"02",X"C2",X"62",X"27",X"3E",X"0F",X"DD",
		X"A6",X"04",X"C2",X"62",X"27",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"AC",X"91",X"FE",X"20",
		X"CA",X"3E",X"2C",X"E6",X"F8",X"FE",X"30",X"CC",X"E3",X"2C",X"3A",X"01",X"48",X"CB",X"7F",X"CA",
		X"62",X"27",X"21",X"00",X"50",X"CB",X"6F",X"28",X"0A",X"3A",X"80",X"50",X"CB",X"47",X"20",X"03",
		X"21",X"40",X"50",X"7E",X"2F",X"E6",X"1F",X"FE",X"10",X"C2",X"62",X"27",X"DD",X"66",X"02",X"DD",
		X"6E",X"04",X"CD",X"AC",X"91",X"FE",X"FF",X"CA",X"62",X"27",X"CB",X"7F",X"C2",X"62",X"27",X"CB",
		X"5F",X"C2",X"62",X"27",X"FD",X"77",X"09",X"E6",X"F0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"FE",X"03",X"20",X"03",X"C3",X"62",X"27",X"CB",X"DE",X"CB",X"FF",X"FD",X"77",X"00",X"FD",
		X"36",X"10",X"00",X"21",X"F1",X"49",X"06",X"08",X"CF",X"21",X"80",X"4A",X"06",X"08",X"CF",X"C3",
		X"62",X"27",X"FD",X"7E",X"01",X"21",X"5B",X"28",X"F7",X"18",X"0A",X"6A",X"28",X"8B",X"28",X"9D",
		X"28",X"8B",X"28",X"9D",X"28",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"04",X"FE",X"41",X"38",
		X"07",X"CD",X"F8",X"2D",X"CD",X"49",X"2E",X"C9",X"FE",X"38",X"30",X"06",X"DD",X"36",X"04",X"FE",
		X"18",X"EF",X"DD",X"7E",X"02",X"FE",X"80",X"28",X"E8",X"18",X"E9",X"3E",X"0F",X"DD",X"A6",X"02",
		X"20",X"15",X"DD",X"7E",X"02",X"FE",X"30",X"38",X"0E",X"FE",X"E1",X"30",X"0A",X"DD",X"36",X"01",
		X"0C",X"FD",X"36",X"01",X"00",X"18",X"C3",X"3E",X"01",X"FD",X"BE",X"01",X"CA",X"CA",X"28",X"C3",
		X"2C",X"29",X"FD",X"7E",X"01",X"21",X"BB",X"28",X"F7",X"18",X"0A",X"EE",X"28",X"CA",X"28",X"EE",
		X"28",X"00",X"29",X"00",X"29",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"02",X"FE",X"E0",X"30",
		X"07",X"CD",X"F8",X"2D",X"CD",X"49",X"2E",X"C9",X"DD",X"7E",X"02",X"FE",X"E2",X"38",X"06",X"DD",
		X"36",X"02",X"22",X"18",X"EC",X"DD",X"7E",X"04",X"FE",X"90",X"28",X"E5",X"18",X"E6",X"3E",X"0F",
		X"DD",X"A6",X"04",X"20",X"15",X"DD",X"7E",X"04",X"FE",X"40",X"38",X"0E",X"FE",X"F1",X"30",X"0A",
		X"DD",X"36",X"01",X"08",X"FD",X"36",X"01",X"01",X"18",X"C0",X"AF",X"FD",X"BE",X"01",X"CA",X"6A",
		X"28",X"C3",X"8E",X"29",X"FD",X"7E",X"01",X"21",X"1D",X"29",X"F7",X"18",X"0A",X"50",X"29",X"62",
		X"29",X"50",X"29",X"2C",X"29",X"62",X"29",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"02",X"FE",
		X"31",X"38",X"07",X"CD",X"F8",X"2D",X"CD",X"49",X"2E",X"C9",X"DD",X"7E",X"02",X"FE",X"28",X"30",
		X"06",X"DD",X"36",X"02",X"EE",X"18",X"EC",X"DD",X"7E",X"04",X"FE",X"90",X"28",X"E5",X"18",X"E6",
		X"3E",X"0F",X"DD",X"A6",X"04",X"20",X"15",X"DD",X"7E",X"04",X"FE",X"40",X"38",X"0E",X"FE",X"F1",
		X"30",X"0A",X"DD",X"36",X"01",X"88",X"FD",X"36",X"01",X"03",X"18",X"C0",X"AF",X"FD",X"BE",X"01",
		X"CA",X"6A",X"28",X"C3",X"8E",X"29",X"FD",X"7E",X"01",X"21",X"7F",X"29",X"F7",X"18",X"0A",X"C1",
		X"29",X"AF",X"29",X"8E",X"29",X"AF",X"29",X"C1",X"29",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",
		X"04",X"FE",X"F8",X"38",X"06",X"DD",X"36",X"04",X"32",X"18",X"04",X"FE",X"F0",X"30",X"07",X"CD",
		X"F8",X"2D",X"CD",X"49",X"2E",X"C9",X"DD",X"7E",X"02",X"FE",X"80",X"28",X"F2",X"18",X"F3",X"3E",
		X"0F",X"DD",X"A6",X"02",X"20",X"15",X"DD",X"7E",X"02",X"FE",X"30",X"38",X"0E",X"FE",X"E1",X"30",
		X"0A",X"DD",X"36",X"01",X"0A",X"FD",X"36",X"01",X"02",X"18",X"C3",X"3E",X"01",X"FD",X"BE",X"01",
		X"CA",X"CA",X"28",X"C3",X"2C",X"29",X"3E",X"0F",X"DD",X"A6",X"02",X"20",X"10",X"3E",X"0F",X"DD",
		X"A6",X"04",X"20",X"09",X"DD",X"36",X"01",X"0E",X"DD",X"36",X"00",X"00",X"C9",X"FD",X"7E",X"01",
		X"DF",X"6A",X"28",X"CA",X"28",X"8E",X"29",X"2C",X"29",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"3E",
		X"FA",X"84",X"57",X"3E",X"06",X"84",X"5F",X"3E",X"FA",X"85",X"67",X"3E",X"06",X"85",X"6F",X"FD",
		X"E5",X"DD",X"E5",X"DD",X"21",X"45",X"48",X"FD",X"21",X"27",X"4A",X"06",X"06",X"0E",X"00",X"DD",
		X"7E",X"02",X"BA",X"38",X"0C",X"BB",X"30",X"09",X"DD",X"7E",X"04",X"BC",X"38",X"03",X"BD",X"38",
		X"18",X"D5",X"11",X"05",X"00",X"DD",X"19",X"3E",X"04",X"B8",X"38",X"05",X"11",X"0E",X"00",X"FD",
		X"19",X"D1",X"10",X"DB",X"DD",X"E1",X"FD",X"E1",X"C9",X"3E",X"04",X"B8",X"38",X"12",X"FD",X"7E",
		X"00",X"FE",X"02",X"CA",X"B5",X"2A",X"FE",X"03",X"28",X"06",X"FE",X"01",X"28",X"02",X"18",X"D1",
		X"DD",X"E1",X"FD",X"E1",X"C1",X"3E",X"80",X"CD",X"40",X"03",X"21",X"A4",X"2C",X"CD",X"91",X"91",
		X"21",X"02",X"48",X"CB",X"6E",X"CB",X"EE",X"3E",X"23",X"06",X"05",X"FF",X"CD",X"82",X"2A",X"C3",
		X"8E",X"2C",X"3E",X"02",X"CD",X"40",X"03",X"21",X"45",X"48",X"06",X"23",X"CF",X"DD",X"36",X"01",
		X"0F",X"DD",X"36",X"00",X"00",X"3E",X"23",X"06",X"28",X"FF",X"DD",X"36",X"01",X"10",X"DD",X"36",
		X"00",X"00",X"3E",X"23",X"06",X"30",X"FF",X"DD",X"36",X"01",X"17",X"DD",X"36",X"00",X"00",X"3E",
		X"23",X"06",X"10",X"FF",X"C9",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"0C",X"CD",X"40",X"03",X"FD",
		X"36",X"00",X"04",X"FD",X"36",X"01",X"40",X"FD",X"36",X"06",X"02",X"FD",X"36",X"04",X"35",X"FD",
		X"21",X"27",X"4A",X"06",X"04",X"FD",X"7E",X"00",X"FE",X"02",X"28",X"11",X"11",X"0E",X"00",X"FD",
		X"19",X"10",X"F2",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"84",X"CD",X"40",X"03",X"21",X"00",X"2B",
		X"CD",X"BA",X"2C",X"C2",X"D5",X"2C",X"DD",X"E1",X"FD",X"E1",X"C9",X"00",X"00",X"00",X"01",X"00",
		X"00",X"FD",X"21",X"F1",X"49",X"FD",X"CB",X"00",X"7E",X"20",X"31",X"CD",X"9A",X"2D",X"28",X"05",
		X"3E",X"04",X"CD",X"40",X"03",X"FD",X"CB",X"00",X"FE",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"E5",
		X"CD",X"AC",X"91",X"CB",X"DE",X"E1",X"CD",X"1E",X"92",X"1E",X"0A",X"3E",X"01",X"01",X"02",X"02",
		X"CD",X"5C",X"90",X"3E",X"16",X"32",X"66",X"48",X"CD",X"A9",X"2E",X"C9",X"FD",X"7E",X"01",X"B7",
		X"28",X"04",X"FD",X"35",X"01",X"C9",X"CD",X"C7",X"2E",X"C0",X"CD",X"9A",X"2D",X"28",X"05",X"3E",
		X"81",X"CD",X"40",X"03",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"AC",X"91",X"CB",X"FE",X"CB",
		X"9E",X"21",X"63",X"48",X"06",X"05",X"CF",X"AF",X"DD",X"36",X"01",X"0E",X"32",X"E0",X"49",X"DD",
		X"66",X"02",X"DD",X"6E",X"04",X"CD",X"6E",X"AF",X"C9",X"FD",X"21",X"F1",X"49",X"FD",X"CB",X"00",
		X"7E",X"20",X"47",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"04",X"CD",X"40",X"03",X"FD",X"CB",X"00",
		X"FE",X"3A",X"E9",X"49",X"E6",X"07",X"5F",X"3A",X"01",X"48",X"CB",X"57",X"7B",X"28",X"05",X"CD",
		X"87",X"95",X"18",X"03",X"CD",X"76",X"95",X"57",X"D5",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"E5",
		X"CD",X"AC",X"91",X"CB",X"DE",X"E1",X"CD",X"1E",X"92",X"D1",X"7A",X"01",X"02",X"02",X"CD",X"5C",
		X"90",X"3E",X"16",X"32",X"66",X"48",X"CD",X"A9",X"2E",X"C9",X"FD",X"7E",X"01",X"B7",X"28",X"04",
		X"FD",X"35",X"01",X"C9",X"CD",X"C7",X"2E",X"C0",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"81",X"CD",
		X"40",X"03",X"21",X"A3",X"49",X"34",X"DD",X"36",X"01",X"0E",X"DD",X"66",X"02",X"DD",X"6E",X"04",
		X"CD",X"AC",X"91",X"CB",X"FE",X"CB",X"9E",X"CD",X"90",X"3F",X"21",X"63",X"48",X"06",X"05",X"CF",
		X"AF",X"32",X"E0",X"49",X"3A",X"E9",X"49",X"E6",X"07",X"3D",X"21",X"18",X"2C",X"CD",X"1D",X"94",
		X"EB",X"CD",X"BA",X"2C",X"C2",X"D5",X"2C",X"C9",X"25",X"2C",X"2B",X"2C",X"31",X"2C",X"37",X"2C",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"21",X"02",
		X"48",X"CB",X"6E",X"CB",X"EE",X"3E",X"80",X"CD",X"40",X"03",X"3E",X"03",X"CD",X"40",X"03",X"21",
		X"A4",X"2C",X"CD",X"91",X"91",X"3E",X"23",X"06",X"01",X"FF",X"21",X"A8",X"2C",X"7E",X"23",X"DD",
		X"77",X"01",X"DD",X"36",X"00",X"00",X"06",X"04",X"C5",X"3E",X"23",X"06",X"04",X"FF",X"C1",X"7E",
		X"23",X"FE",X"FF",X"20",X"10",X"05",X"28",X"16",X"21",X"A8",X"2C",X"78",X"FE",X"03",X"30",X"EF",
		X"21",X"B1",X"2C",X"18",X"EA",X"DD",X"77",X"01",X"DD",X"36",X"00",X"00",X"18",X"DA",X"DD",X"36",
		X"01",X"00",X"DD",X"36",X"00",X"00",X"3E",X"23",X"06",X"20",X"FF",X"3E",X"00",X"01",X"B8",X"32",
		X"FF",X"3E",X"60",X"FF",X"15",X"16",X"17",X"FF",X"11",X"12",X"13",X"52",X"51",X"D2",X"93",X"92",
		X"FF",X"14",X"15",X"16",X"55",X"54",X"95",X"96",X"D5",X"FF",X"DD",X"E5",X"CD",X"92",X"90",X"DD",
		X"E1",X"21",X"CF",X"2C",X"11",X"88",X"49",X"06",X"06",X"CD",X"80",X"90",X"FE",X"01",X"C9",X"00",
		X"01",X"00",X"00",X"00",X"00",X"3E",X"80",X"CD",X"40",X"03",X"3E",X"00",X"01",X"9F",X"31",X"FF",
		X"3E",X"60",X"FF",X"FD",X"CB",X"0A",X"76",X"C0",X"CD",X"D6",X"0C",X"3A",X"A5",X"49",X"3C",X"32",
		X"A5",X"49",X"FE",X"04",X"28",X"05",X"CD",X"B6",X"2D",X"18",X"18",X"21",X"CE",X"41",X"01",X"02",
		X"02",X"1E",X"16",X"AF",X"CD",X"0C",X"90",X"3A",X"AA",X"48",X"CB",X"7F",X"20",X"05",X"E6",X"07",
		X"32",X"AA",X"48",X"FD",X"E5",X"FD",X"21",X"27",X"4A",X"06",X"04",X"0E",X"00",X"FD",X"7E",X"00",
		X"FE",X"03",X"28",X"04",X"FE",X"02",X"20",X"0C",X"FD",X"36",X"00",X"02",X"CD",X"0E",X"8E",X"CD",
		X"FE",X"88",X"0E",X"01",X"11",X"0E",X"00",X"FD",X"19",X"10",X"E2",X"AF",X"B9",X"28",X"19",X"21",
		X"86",X"2D",X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"CD",X"1D",X"94",X"ED",
		X"53",X"25",X"4A",X"3E",X"15",X"CD",X"40",X"03",X"FD",X"E1",X"21",X"7C",X"2D",X"3A",X"AA",X"49",
		X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"CB",X"0A",X"F6",
		X"FD",X"77",X"0F",X"FD",X"36",X"02",X"FF",X"FD",X"36",X"03",X"FF",X"C9",X"2D",X"2D",X"2D",X"2D",
		X"2D",X"2D",X"2D",X"2D",X"2D",X"2D",X"69",X"01",X"2D",X"01",X"2D",X"01",X"69",X"01",X"2D",X"01",
		X"F0",X"00",X"2D",X"01",X"F0",X"00",X"B4",X"00",X"B4",X"00",X"2A",X"25",X"48",X"11",X"D9",X"A3",
		X"B7",X"E5",X"ED",X"52",X"E1",X"C8",X"11",X"BD",X"A4",X"B7",X"E5",X"ED",X"52",X"E1",X"C8",X"11",
		X"FB",X"9E",X"B7",X"ED",X"52",X"C9",X"3A",X"A5",X"49",X"FE",X"04",X"D0",X"21",X"CE",X"2D",X"CD",
		X"1D",X"94",X"7B",X"5A",X"21",X"CE",X"41",X"01",X"02",X"02",X"CD",X"5C",X"90",X"C9",X"60",X"18",
		X"64",X"0C",X"68",X"15",X"6C",X"15",X"21",X"EE",X"2D",X"3A",X"AA",X"49",X"FE",X"05",X"38",X"02",
		X"3E",X"05",X"3D",X"CD",X"17",X"94",X"5E",X"23",X"56",X"EB",X"22",X"E2",X"49",X"C9",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FD",X"7E",X"0E",X"CB",X"BF",X"B7",X"20",X"22",
		X"3E",X"02",X"FD",X"B6",X"0E",X"FD",X"77",X"0E",X"3E",X"10",X"FD",X"CB",X"0E",X"7E",X"FD",X"CB",
		X"0E",X"FE",X"28",X"06",X"3E",X"01",X"FD",X"CB",X"0E",X"BE",X"CD",X"9A",X"2D",X"28",X"03",X"CD",
		X"40",X"03",X"FD",X"35",X"0E",X"21",X"41",X"2E",X"FD",X"7E",X"01",X"CD",X"17",X"94",X"4E",X"23",
		X"46",X"DD",X"66",X"02",X"DD",X"6E",X"04",X"CD",X"A5",X"91",X"DD",X"74",X"02",X"DD",X"75",X"04",
		X"C9",X"00",X"FE",X"02",X"00",X"00",X"02",X"FE",X"00",X"21",X"5E",X"2E",X"FD",X"7E",X"01",X"CD",
		X"17",X"94",X"DD",X"7E",X"01",X"BE",X"20",X"01",X"23",X"7E",X"DD",X"77",X"01",X"C9",X"0C",X"0D",
		X"08",X"09",X"0A",X"0B",X"88",X"89",X"3A",X"01",X"48",X"CB",X"7F",X"28",X"16",X"CB",X"6F",X"21",
		X"00",X"50",X"28",X"0A",X"3A",X"80",X"50",X"CB",X"47",X"20",X"03",X"21",X"40",X"50",X"7E",X"2F",
		X"E6",X"0F",X"C9",X"3A",X"E0",X"4A",X"B7",X"20",X"13",X"2A",X"E2",X"4A",X"23",X"22",X"E2",X"4A",
		X"7E",X"B7",X"CA",X"A5",X"2E",X"32",X"E0",X"4A",X"23",X"22",X"E2",X"4A",X"21",X"E0",X"4A",X"35",
		X"2A",X"E2",X"4A",X"7E",X"C9",X"C1",X"CA",X"0C",X"28",X"DD",X"7E",X"02",X"32",X"65",X"48",X"DD",
		X"7E",X"04",X"32",X"67",X"48",X"3E",X"18",X"32",X"64",X"48",X"AF",X"32",X"63",X"48",X"DD",X"36",
		X"01",X"01",X"FD",X"36",X"01",X"01",X"C9",X"FD",X"36",X"01",X"01",X"DD",X"34",X"01",X"3A",X"64",
		X"48",X"3C",X"32",X"64",X"48",X"F5",X"AF",X"32",X"63",X"48",X"F1",X"FE",X"1F",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"18",X"06",X"31",X"C0",X"4F",X"C3",X"32",X"2F",X"31",X"C0",X"4F",X"CD",X"D5",X"04",X"CD",X"40",
		X"36",X"79",X"32",X"04",X"48",X"21",X"DD",X"38",X"11",X"00",X"4C",X"01",X"F0",X"00",X"ED",X"B0",
		X"21",X"DD",X"38",X"11",X"08",X"48",X"01",X"06",X"00",X"ED",X"B0",X"EF",X"CD",X"CB",X"34",X"21",
		X"E8",X"36",X"CD",X"91",X"91",X"AF",X"32",X"01",X"48",X"CD",X"14",X"36",X"CD",X"43",X"35",X"CD",
		X"80",X"3A",X"CD",X"CB",X"34",X"21",X"01",X"48",X"7E",X"E6",X"80",X"77",X"23",X"36",X"00",X"CD",
		X"14",X"36",X"21",X"E8",X"36",X"CD",X"91",X"91",X"CD",X"43",X"35",X"CD",X"DC",X"35",X"CD",X"6F",
		X"35",X"3A",X"01",X"48",X"CB",X"7F",X"CA",X"90",X"30",X"FD",X"21",X"05",X"48",X"FD",X"7E",X"00",
		X"B7",X"20",X"0D",X"E7",X"21",X"01",X"48",X"36",X"00",X"23",X"36",X"00",X"EF",X"C3",X"1C",X"2F",
		X"DD",X"21",X"5A",X"37",X"CD",X"0A",X"8F",X"21",X"49",X"42",X"DD",X"21",X"06",X"48",X"1E",X"02",
		X"06",X"02",X"0E",X"FF",X"CD",X"1E",X"90",X"DD",X"21",X"01",X"38",X"CD",X"0A",X"8F",X"DD",X"21",
		X"18",X"38",X"CD",X"0A",X"8F",X"CD",X"40",X"36",X"FE",X"06",X"CA",X"FA",X"2F",X"DD",X"21",X"D2",
		X"37",X"CD",X"0A",X"8F",X"FD",X"7E",X"00",X"FE",X"01",X"20",X"24",X"DD",X"21",X"8B",X"37",X"CD",
		X"0A",X"8F",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"40",X"50",X"CB",X"6F",X"20",X"E6",X"FD",X"35",
		X"00",X"21",X"E3",X"36",X"11",X"07",X"48",X"06",X"02",X"CD",X"EF",X"8F",X"C3",X"74",X"30",X"DD",
		X"21",X"A1",X"37",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"40",X"50",X"CB",X"6F",
		X"28",X"DC",X"CB",X"77",X"20",X"F0",X"FD",X"35",X"00",X"FD",X"35",X"00",X"21",X"E5",X"36",X"11",
		X"07",X"48",X"06",X"02",X"CD",X"EF",X"8F",X"C3",X"6D",X"30",X"FD",X"7E",X"00",X"FE",X"02",X"30",
		X"0E",X"DD",X"21",X"C2",X"37",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"01",X"FF",X"18",X"EB",X"DD",
		X"21",X"D2",X"37",X"CD",X"0A",X"8F",X"FD",X"7E",X"00",X"FE",X"04",X"30",X"26",X"DD",X"21",X"8B",
		X"37",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"40",X"50",X"CB",X"6F",X"20",X"E6",
		X"FD",X"35",X"00",X"FD",X"35",X"00",X"21",X"E5",X"36",X"11",X"07",X"48",X"06",X"02",X"CD",X"EF",
		X"8F",X"18",X"31",X"DD",X"21",X"A1",X"37",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"01",X"FF",X"3A",
		X"40",X"50",X"CB",X"6F",X"28",X"DA",X"CB",X"77",X"20",X"F0",X"FD",X"7E",X"00",X"D6",X"04",X"FD",
		X"77",X"00",X"21",X"E7",X"36",X"11",X"07",X"48",X"06",X"02",X"CD",X"EF",X"8F",X"21",X"01",X"48",
		X"CB",X"76",X"CB",X"F6",X"21",X"02",X"48",X"CB",X"7E",X"CB",X"FE",X"21",X"49",X"42",X"DD",X"21",
		X"06",X"48",X"1E",X"02",X"06",X"02",X"0E",X"FF",X"CD",X"1E",X"90",X"3E",X"23",X"06",X"04",X"FF",
		X"3A",X"01",X"48",X"CB",X"7F",X"28",X"06",X"21",X"0E",X"48",X"06",X"0C",X"CF",X"21",X"0B",X"37",
		X"11",X"88",X"49",X"01",X"24",X"00",X"ED",X"B0",X"21",X"0B",X"37",X"11",X"B0",X"49",X"01",X"24",
		X"00",X"ED",X"B0",X"3A",X"80",X"50",X"2F",X"E6",X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"C6",X"03",X"32",X"A7",X"49",X"32",X"CF",X"49",X"CD",X"36",X"92",X"21",X"68",X"48",X"11",
		X"F8",X"48",X"01",X"90",X"00",X"ED",X"B0",X"CD",X"36",X"92",X"21",X"68",X"48",X"11",X"68",X"48",
		X"FD",X"21",X"D0",X"4A",X"CD",X"9A",X"36",X"21",X"F8",X"48",X"11",X"F8",X"48",X"FD",X"21",X"F0",
		X"4A",X"CD",X"9A",X"36",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"16",X"21",X"41",X"38",X"11",X"68",
		X"48",X"01",X"90",X"00",X"ED",X"B0",X"11",X"D0",X"4A",X"21",X"D1",X"38",X"01",X"0C",X"00",X"ED",
		X"B0",X"CD",X"14",X"36",X"CD",X"43",X"35",X"CD",X"CB",X"34",X"CD",X"DC",X"35",X"CD",X"6F",X"35",
		X"CD",X"F0",X"14",X"3E",X"23",X"06",X"40",X"FF",X"CD",X"5B",X"35",X"CD",X"CE",X"34",X"CD",X"5F",
		X"36",X"3A",X"A4",X"49",X"B7",X"28",X"0D",X"CD",X"2D",X"95",X"CD",X"CE",X"34",X"3E",X"23",X"06",
		X"40",X"FF",X"18",X"12",X"3E",X"12",X"CD",X"40",X"03",X"CD",X"D7",X"94",X"3E",X"23",X"06",X"08",
		X"FF",X"3E",X"80",X"CD",X"40",X"03",X"CD",X"5B",X"35",X"CD",X"5F",X"36",X"CD",X"3D",X"94",X"21",
		X"F1",X"36",X"CD",X"99",X"91",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"03",X"3E",X"60",X"FF",X"DD",
		X"21",X"67",X"37",X"21",X"70",X"37",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"07",X"DD",X"21",X"79",
		X"37",X"21",X"82",X"37",X"DD",X"E5",X"E5",X"E5",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"18",X"FF",
		X"DD",X"E1",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"10",X"FF",X"E1",X"DD",X"E1",X"18",X"E5",X"31",
		X"C0",X"4F",X"21",X"E8",X"36",X"CD",X"91",X"91",X"3E",X"80",X"CD",X"40",X"03",X"3E",X"16",X"CD",
		X"40",X"03",X"DD",X"21",X"67",X"37",X"3A",X"01",X"48",X"CB",X"6F",X"28",X"04",X"DD",X"21",X"79",
		X"37",X"CD",X"0A",X"8F",X"21",X"02",X"48",X"7E",X"E6",X"80",X"77",X"2B",X"7E",X"E6",X"F8",X"77",
		X"3E",X"01",X"01",X"00",X"3A",X"FF",X"3E",X"23",X"06",X"20",X"FF",X"21",X"40",X"48",X"06",X"28",
		X"CF",X"CD",X"2D",X"95",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"2C",X"48",X"CB",X"7F",X"20",X"F4",
		X"3E",X"23",X"06",X"20",X"FF",X"CD",X"06",X"34",X"3A",X"AA",X"49",X"3C",X"20",X"02",X"3E",X"01",
		X"32",X"AA",X"49",X"21",X"88",X"49",X"06",X"06",X"CF",X"CD",X"6F",X"35",X"3E",X"11",X"FF",X"CD",
		X"5B",X"35",X"CD",X"CB",X"34",X"21",X"07",X"37",X"CD",X"99",X"91",X"3E",X"30",X"FF",X"3E",X"80",
		X"FF",X"F5",X"FE",X"10",X"28",X"06",X"21",X"88",X"49",X"06",X"06",X"CF",X"3A",X"01",X"48",X"CB",
		X"7F",X"20",X"25",X"3E",X"23",X"06",X"40",X"FF",X"CD",X"43",X"35",X"CD",X"80",X"A5",X"3E",X"23",
		X"06",X"3C",X"FF",X"DD",X"21",X"01",X"38",X"CD",X"0A",X"8F",X"3E",X"23",X"06",X"C0",X"FF",X"C3",
		X"1C",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"CD",X"6D",X"34",X"21",X"B1",X"32",X"11",X"A9",
		X"49",X"06",X"02",X"CD",X"DA",X"8F",X"21",X"0B",X"37",X"11",X"88",X"49",X"01",X"1E",X"00",X"ED",
		X"B0",X"3A",X"A6",X"49",X"E6",X"0F",X"32",X"A6",X"49",X"CD",X"36",X"92",X"21",X"68",X"48",X"11",
		X"68",X"48",X"FD",X"21",X"D0",X"4A",X"CD",X"9A",X"36",X"F1",X"FE",X"20",X"20",X"1A",X"3A",X"A7",
		X"49",X"FE",X"02",X"30",X"0B",X"21",X"B1",X"32",X"11",X"A9",X"49",X"06",X"02",X"CD",X"EF",X"8F",
		X"3E",X"23",X"06",X"40",X"FF",X"C3",X"F9",X"32",X"3E",X"23",X"06",X"80",X"FF",X"C3",X"11",X"31",
		X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"31",X"C0",X"4F",X"21",X"E8",X"36",X"CD",X"91",
		X"91",X"3E",X"80",X"CD",X"40",X"03",X"DD",X"21",X"67",X"37",X"3A",X"01",X"48",X"CB",X"6F",X"28",
		X"04",X"DD",X"21",X"79",X"37",X"CD",X"0A",X"8F",X"21",X"02",X"48",X"7E",X"E6",X"80",X"77",X"2B",
		X"7E",X"E6",X"F8",X"77",X"3E",X"23",X"06",X"30",X"FF",X"3A",X"01",X"48",X"CB",X"7F",X"CA",X"03",
		X"32",X"21",X"A4",X"49",X"34",X"AF",X"32",X"96",X"49",X"11",X"01",X"48",X"1A",X"E6",X"F8",X"12",
		X"21",X"A7",X"49",X"1A",X"CB",X"77",X"20",X"18",X"35",X"C2",X"11",X"31",X"CD",X"14",X"35",X"CD",
		X"C1",X"33",X"3E",X"23",X"06",X"20",X"FF",X"CD",X"43",X"35",X"CD",X"10",X"17",X"C3",X"32",X"2F",
		X"35",X"21",X"CF",X"49",X"28",X"07",X"7E",X"B7",X"CA",X"11",X"31",X"18",X"1A",X"CD",X"14",X"35",
		X"CD",X"C1",X"33",X"3E",X"23",X"06",X"20",X"FF",X"CD",X"43",X"35",X"CD",X"10",X"17",X"3A",X"CF",
		X"49",X"B7",X"20",X"03",X"C3",X"32",X"2F",X"3A",X"01",X"48",X"CB",X"6F",X"CB",X"EF",X"28",X"02",
		X"CB",X"AF",X"32",X"01",X"48",X"21",X"88",X"49",X"11",X"E0",X"49",X"01",X"24",X"00",X"ED",X"B0",
		X"21",X"B0",X"49",X"11",X"88",X"49",X"01",X"24",X"00",X"ED",X"B0",X"21",X"E0",X"49",X"11",X"B0",
		X"49",X"01",X"24",X"00",X"ED",X"B0",X"21",X"D0",X"4A",X"11",X"E0",X"49",X"01",X"10",X"00",X"ED",
		X"B0",X"21",X"F0",X"4A",X"11",X"D0",X"4A",X"01",X"10",X"00",X"ED",X"B0",X"21",X"E0",X"49",X"11",
		X"F0",X"4A",X"01",X"10",X"00",X"ED",X"B0",X"21",X"68",X"48",X"11",X"E0",X"49",X"01",X"90",X"00",
		X"ED",X"B0",X"21",X"F8",X"48",X"11",X"68",X"48",X"01",X"90",X"00",X"ED",X"B0",X"21",X"E0",X"49",
		X"11",X"F8",X"48",X"01",X"90",X"00",X"ED",X"B0",X"21",X"E0",X"49",X"06",X"90",X"CF",X"C3",X"11",
		X"31",X"21",X"0E",X"48",X"11",X"14",X"48",X"06",X"06",X"CD",X"80",X"90",X"21",X"0E",X"48",X"FE",
		X"02",X"38",X"03",X"21",X"14",X"48",X"E5",X"11",X"08",X"48",X"06",X"06",X"CD",X"80",X"90",X"E1",
		X"FE",X"01",X"20",X"08",X"11",X"08",X"48",X"01",X"06",X"00",X"ED",X"B0",X"21",X"DF",X"41",X"DD",
		X"21",X"08",X"48",X"1E",X"17",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",X"88",X"49",X"06",
		X"06",X"CF",X"CD",X"6F",X"35",X"C9",X"3E",X"1D",X"CD",X"40",X"03",X"21",X"B2",X"32",X"11",X"8E",
		X"49",X"06",X"06",X"CD",X"80",X"90",X"FE",X"02",X"20",X"2A",X"21",X"B7",X"32",X"CD",X"92",X"90",
		X"21",X"B7",X"32",X"11",X"93",X"49",X"06",X"06",X"CD",X"EF",X"8F",X"3A",X"FC",X"46",X"5F",X"21",
		X"FC",X"42",X"DD",X"21",X"8E",X"49",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"3E",X"23",X"06",
		X"02",X"FF",X"18",X"C7",X"3E",X"81",X"CD",X"40",X"03",X"21",X"93",X"49",X"CD",X"92",X"90",X"21",
		X"8E",X"49",X"06",X"06",X"CF",X"3A",X"FC",X"46",X"5F",X"21",X"FC",X"42",X"DD",X"21",X"8E",X"49",
		X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"3E",X"23",X"06",X"40",X"FF",X"C9",X"3E",X"1D",X"CD",
		X"40",X"03",X"21",X"B2",X"32",X"11",X"88",X"49",X"06",X"06",X"CD",X"80",X"90",X"FE",X"02",X"20",
		X"28",X"21",X"B7",X"32",X"CD",X"AC",X"90",X"21",X"B7",X"32",X"11",X"8D",X"49",X"06",X"06",X"CD",
		X"EF",X"8F",X"21",X"BD",X"41",X"DD",X"21",X"88",X"49",X"1E",X"04",X"06",X"06",X"0E",X"00",X"CD",
		X"1E",X"90",X"3E",X"23",X"06",X"02",X"FF",X"18",X"C9",X"3E",X"81",X"CD",X"40",X"03",X"21",X"8D",
		X"49",X"CD",X"AC",X"90",X"21",X"88",X"49",X"06",X"06",X"CF",X"21",X"BD",X"41",X"DD",X"21",X"88",
		X"49",X"1E",X"04",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"C9",X"AF",X"18",X"2A",X"3A",X"AA",
		X"49",X"FE",X"09",X"38",X"04",X"D6",X"08",X"18",X"F8",X"0E",X"00",X"FE",X"03",X"38",X"05",X"0C",
		X"D6",X"02",X"18",X"F7",X"79",X"81",X"4F",X"06",X"00",X"21",X"FF",X"34",X"09",X"7E",X"23",X"32",
		X"05",X"50",X"7E",X"32",X"06",X"50",X"3E",X"01",X"21",X"01",X"50",X"77",X"23",X"77",X"C9",X"01",
		X"00",X"00",X"01",X"01",X"01",X"00",X"00",X"11",X"13",X"48",X"3A",X"01",X"48",X"CB",X"6F",X"C8",
		X"11",X"19",X"48",X"C9",X"E5",X"D5",X"21",X"CE",X"40",X"01",X"14",X"03",X"AF",X"1E",X"00",X"CD",
		X"4A",X"90",X"21",X"EF",X"40",X"06",X"12",X"1E",X"00",X"DD",X"21",X"DD",X"37",X"3A",X"01",X"48",
		X"CB",X"6F",X"28",X"04",X"DD",X"21",X"EF",X"37",X"CD",X"7D",X"8F",X"D1",X"E1",X"3E",X"23",X"06",
		X"40",X"FF",X"C9",X"21",X"00",X"40",X"01",X"00",X"04",X"1E",X"00",X"CD",X"02",X"8F",X"21",X"00",
		X"44",X"01",X"00",X"04",X"1E",X"00",X"CD",X"02",X"8F",X"18",X"0D",X"21",X"00",X"40",X"01",X"20",
		X"1C",X"1E",X"00",X"3E",X"00",X"CD",X"0C",X"90",X"21",X"40",X"48",X"06",X"28",X"CF",X"C9",X"21",
		X"BF",X"40",X"DD",X"21",X"0E",X"48",X"1E",X"05",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",
		X"FF",X"42",X"DD",X"21",X"14",X"48",X"1E",X"05",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",
		X"BD",X"41",X"DD",X"21",X"88",X"49",X"1E",X"04",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",
		X"DF",X"41",X"DD",X"21",X"08",X"48",X"1E",X"17",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"21",
		X"FD",X"40",X"DD",X"21",X"A8",X"49",X"1E",X"02",X"06",X"02",X"0E",X"00",X"CD",X"1E",X"90",X"CD",
		X"FC",X"35",X"3A",X"A6",X"49",X"CB",X"67",X"1E",X"05",X"28",X"02",X"1E",X"02",X"21",X"FC",X"42",
		X"DD",X"21",X"8E",X"49",X"06",X"06",X"0E",X"00",X"CD",X"1E",X"90",X"C9",X"DD",X"21",X"2F",X"37",
		X"CD",X"0A",X"8F",X"21",X"5C",X"41",X"01",X"0C",X"03",X"3E",X"51",X"1E",X"10",X"CD",X"4A",X"90",
		X"21",X"7D",X"41",X"01",X"0A",X"01",X"AF",X"5F",X"CD",X"0C",X"90",X"C9",X"3A",X"A7",X"49",X"B7",
		X"C8",X"47",X"3A",X"A4",X"49",X"B7",X"20",X"07",X"3A",X"AA",X"49",X"FE",X"02",X"38",X"01",X"05",
		X"CD",X"70",X"91",X"C9",X"21",X"01",X"48",X"3A",X"80",X"50",X"2F",X"E6",X"03",X"CB",X"6E",X"28",
		X"02",X"CB",X"D7",X"21",X"32",X"36",X"06",X"00",X"4F",X"09",X"7E",X"32",X"03",X"50",X"32",X"1B",
		X"48",X"C9",X"00",X"00",X"01",X"01",X"00",X"01",X"01",X"00",X"3A",X"01",X"48",X"CB",X"6F",X"C9",
		X"3A",X"80",X"50",X"2F",X"CB",X"07",X"CB",X"07",X"CB",X"07",X"E6",X"06",X"4F",X"21",X"57",X"36",
		X"06",X"00",X"09",X"46",X"23",X"4E",X"C9",X"01",X"01",X"01",X"02",X"01",X"03",X"02",X"01",X"21",
		X"40",X"40",X"DD",X"21",X"10",X"07",X"1E",X"02",X"CD",X"8C",X"8F",X"21",X"4E",X"40",X"1E",X"03",
		X"01",X"02",X"02",X"3E",X"98",X"CD",X"5C",X"90",X"21",X"8E",X"43",X"01",X"02",X"02",X"3E",X"94",
		X"CD",X"5C",X"90",X"21",X"C0",X"41",X"01",X"02",X"02",X"3E",X"9C",X"CD",X"5C",X"90",X"21",X"DA",
		X"41",X"01",X"02",X"02",X"3E",X"90",X"CD",X"5C",X"90",X"C9",X"06",X"90",X"C5",X"7E",X"E6",X"70",
		X"FE",X"10",X"28",X"05",X"23",X"C1",X"10",X"F4",X"C9",X"E5",X"B7",X"ED",X"52",X"7D",X"D5",X"CD",
		X"EA",X"91",X"D1",X"ED",X"5F",X"E6",X"03",X"4F",X"CB",X"47",X"28",X"10",X"06",X"03",X"7C",X"FE",
		X"C0",X"30",X"17",X"06",X"01",X"FE",X"60",X"38",X"11",X"41",X"18",X"0E",X"06",X"00",X"7D",X"FE",
		X"D0",X"30",X"07",X"06",X"02",X"FE",X"60",X"38",X"01",X"41",X"FD",X"70",X"00",X"FD",X"23",X"E1",
		X"18",X"C2",X"00",X"01",X"00",X"02",X"00",X"04",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",
		X"FF",X"02",X"00",X"A5",X"01",X"00",X"AD",X"04",X"A0",X"26",X"06",X"00",X"80",X"05",X"00",X"86",
		X"07",X"20",X"0D",X"08",X"40",X"3F",X"FF",X"01",X"A0",X"18",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",
		X"02",X"7F",X"40",X"00",X"00",X"31",X"50",X"02",X"BF",X"42",X"00",X"00",X"32",X"50",X"02",X"9F",
		X"41",X"00",X"00",X"48",X"49",X"05",X"5D",X"40",X"00",X"00",X"52",X"4F",X"55",X"4E",X"44",X"05",
		X"1D",X"43",X"00",X"00",X"42",X"4F",X"4E",X"55",X"53",X"00",X"00",X"06",X"69",X"41",X"00",X"00",
		X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"00",X"02",X"7F",X"40",X"00",X"00",X"31",X"50",X"00",
		X"00",X"02",X"7F",X"40",X"00",X"00",X"20",X"20",X"00",X"00",X"02",X"BF",X"42",X"00",X"00",X"32",
		X"50",X"00",X"00",X"02",X"BF",X"42",X"00",X"00",X"20",X"20",X"00",X"00",X"0F",X"2F",X"41",X"00",
		X"00",X"31",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"00",X"00",X"0F",X"2F",X"41",X"00",X"00",X"31",X"20",X"4F",X"52",X"20",X"32",X"20",X"50",X"4C",
		X"41",X"59",X"45",X"52",X"53",X"20",X"06",X"AD",X"41",X"00",X"05",X"42",X"55",X"54",X"54",X"4F",
		X"4E",X"00",X"00",X"09",X"6F",X"41",X"00",X"00",X"4D",X"4F",X"52",X"45",X"20",X"43",X"4F",X"49",
		X"4E",X"00",X"00",X"04",X"D1",X"41",X"00",X"05",X"50",X"55",X"53",X"48",X"00",X"47",X"41",X"4D",
		X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"3B",X"31",X"47",
		X"41",X"4D",X"45",X"20",X"4F",X"56",X"45",X"52",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"3B",
		X"32",X"00",X"10",X"01",X"41",X"00",X"17",X"40",X"20",X"31",X"39",X"38",X"32",X"20",X"53",X"41",
		X"4E",X"52",X"49",X"54",X"53",X"55",X"20",X"00",X"00",X"04",X"D7",X"41",X"00",X"00",X"50",X"4C",
		X"41",X"59",X"0D",X"55",X"41",X"01",X"02",X"44",X"14",X"52",X"03",X"45",X"04",X"41",X"05",X"4D",
		X"00",X"3B",X"05",X"53",X"05",X"48",X"05",X"4F",X"05",X"50",X"05",X"50",X"05",X"45",X"05",X"52",
		X"00",X"01",X"02",X"04",X"02",X"03",X"04",X"02",X"03",X"02",X"03",X"04",X"01",X"04",X"02",X"12",
		X"04",X"01",X"01",X"01",X"04",X"13",X"02",X"03",X"04",X"02",X"04",X"03",X"03",X"04",X"02",X"20",
		X"01",X"03",X"04",X"04",X"03",X"03",X"14",X"02",X"04",X"03",X"40",X"04",X"03",X"14",X"01",X"03",
		X"12",X"04",X"02",X"03",X"11",X"04",X"03",X"02",X"04",X"04",X"04",X"02",X"04",X"01",X"04",X"20",
		X"03",X"04",X"02",X"31",X"04",X"02",X"20",X"04",X"03",X"04",X"02",X"03",X"04",X"01",X"02",X"04",
		X"02",X"03",X"03",X"04",X"01",X"13",X"03",X"03",X"02",X"03",X"04",X"02",X"03",X"40",X"04",X"02",
		X"03",X"04",X"02",X"04",X"03",X"40",X"02",X"04",X"11",X"02",X"03",X"04",X"14",X"01",X"04",X"02",
		X"03",X"04",X"02",X"20",X"03",X"04",X"01",X"03",X"04",X"04",X"03",X"11",X"04",X"01",X"04",X"13",
		X"04",X"03",X"04",X"12",X"04",X"02",X"04",X"03",X"02",X"03",X"04",X"03",X"01",X"02",X"03",X"03",
		X"02",X"00",X"01",X"00",X"02",X"02",X"00",X"00",X"03",X"02",X"03",X"03",X"02",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"08",X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"07",
		X"05",X"00",X"00",X"00",X"03",X"00",X"02",X"05",X"04",X"00",X"00",X"00",X"03",X"00",X"02",X"04",
		X"08",X"06",X"00",X"00",X"03",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"03",X"00",X"02",X"01",
		X"01",X"02",X"00",X"00",X"02",X"00",X"02",X"00",X"05",X"06",X"00",X"00",X"02",X"00",X"01",X"09",
		X"08",X"08",X"00",X"00",X"02",X"00",X"01",X"09",X"08",X"00",X"00",X"00",X"02",X"00",X"01",X"08",
		X"05",X"07",X"00",X"00",X"02",X"00",X"01",X"06",X"06",X"03",X"00",X"00",X"02",X"00",X"01",X"05",
		X"00",X"00",X"00",X"00",X"02",X"00",X"01",X"04",X"09",X"09",X"00",X"00",X"02",X"00",X"01",X"03",
		X"05",X"00",X"00",X"00",X"02",X"00",X"01",X"02",X"02",X"02",X"00",X"00",X"02",X"00",X"01",X"01",
		X"05",X"09",X"00",X"00",X"02",X"00",X"01",X"00",X"04",X"02",X"00",X"00",X"02",X"00",X"00",X"09",
		X"09",X"00",X"00",X"00",X"01",X"00",X"00",X"09",X"07",X"05",X"00",X"00",X"01",X"00",X"00",X"09",
		X"05",X"00",X"00",X"00",X"01",X"00",X"00",X"09",X"01",X"05",X"00",X"00",X"01",X"00",X"00",X"08",
		X"07",X"00",X"00",X"00",X"01",X"00",X"00",X"07",X"05",X"00",X"00",X"00",X"01",X"00",X"00",X"07",
		X"06",X"05",X"00",X"00",X"01",X"00",X"00",X"07",X"03",X"00",X"00",X"00",X"01",X"00",X"00",X"06",
		X"00",X"05",X"00",X"00",X"01",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"05",
		X"08",X"00",X"00",X"00",X"01",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"01",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"60",X"4F",X"0E",X"0D",X"CD",X"20",X"3A",X"1E",X"10",X"3E",X"23",X"06",X"02",X"FF",X"4B",
		X"D5",X"CD",X"20",X"3A",X"D1",X"7B",X"3D",X"5F",X"FE",X"0C",X"20",X"EE",X"1E",X"10",X"18",X"EA",
		X"06",X"04",X"21",X"68",X"3A",X"C5",X"79",X"4E",X"23",X"46",X"23",X"5E",X"23",X"56",X"23",X"E5",
		X"C5",X"E1",X"4F",X"CD",X"3B",X"3A",X"E1",X"C1",X"10",X"EB",X"C9",X"06",X"1A",X"7E",X"FE",X"03",
		X"28",X"0F",X"71",X"E5",X"D5",X"16",X"00",X"CB",X"7B",X"28",X"02",X"16",X"FF",X"19",X"71",X"D1",
		X"E1",X"D5",X"5A",X"16",X"00",X"CB",X"7B",X"28",X"02",X"16",X"FF",X"19",X"D1",X"0C",X"79",X"FE",
		X"11",X"20",X"02",X"0E",X"0D",X"10",X"D6",X"C9",X"5A",X"44",X"01",X"20",X"9B",X"47",X"20",X"FF",
		X"A1",X"47",X"FF",X"E0",X"40",X"44",X"20",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FD",X"21",X"37",X"3D",X"FD",X"6E",X"00",X"FD",X"23",X"FD",X"66",X"00",X"FD",X"23",X"FD",X"4E",
		X"00",X"FD",X"23",X"FD",X"7E",X"00",X"FD",X"23",X"5F",X"E6",X"0F",X"47",X"7B",X"E6",X"F0",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"E5",X"21",X"D7",X"3A",X"CD",X"1D",X"94",X"E1",X"19",
		X"FD",X"7E",X"00",X"FD",X"23",X"77",X"CB",X"D4",X"71",X"CB",X"94",X"C5",X"3E",X"23",X"06",X"02",
		X"FF",X"C1",X"10",X"EB",X"FD",X"7E",X"00",X"FE",X"FF",X"28",X"14",X"FE",X"80",X"28",X"04",X"FD",
		X"23",X"18",X"C0",X"FD",X"23",X"18",X"AD",X"01",X"00",X"20",X"00",X"FF",X"FF",X"E0",X"FF",X"3E",
		X"51",X"1E",X"10",X"01",X"01",X"07",X"21",X"72",X"40",X"CD",X"4A",X"90",X"21",X"92",X"40",X"11",
		X"98",X"40",X"0E",X"10",X"06",X"18",X"3E",X"51",X"C5",X"06",X"02",X"77",X"CB",X"D4",X"71",X"CB",
		X"94",X"CD",X"79",X"90",X"EB",X"10",X"F4",X"3E",X"23",X"06",X"02",X"FF",X"C1",X"10",X"E7",X"21",
		X"92",X"43",X"1E",X"10",X"3E",X"51",X"01",X"01",X"07",X"CD",X"4A",X"90",X"21",X"00",X"4B",X"06",
		X"0C",X"CF",X"21",X"E0",X"49",X"06",X"20",X"CF",X"FD",X"21",X"E0",X"49",X"DD",X"21",X"40",X"48",
		X"DD",X"36",X"01",X"0E",X"DD",X"36",X"02",X"10",X"DD",X"36",X"03",X"81",X"DD",X"36",X"04",X"F0",
		X"DD",X"36",X"00",X"00",X"FD",X"36",X"02",X"88",X"FD",X"36",X"03",X"88",X"11",X"D3",X"45",X"ED",
		X"53",X"05",X"4B",X"21",X"13",X"46",X"22",X"03",X"4B",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",
		X"E0",X"49",X"DD",X"21",X"40",X"48",X"FD",X"7E",X"00",X"FE",X"01",X"28",X"26",X"3E",X"80",X"DD",
		X"BE",X"02",X"20",X"11",X"DD",X"36",X"01",X"0E",X"DD",X"36",X"00",X"00",X"FD",X"34",X"00",X"FD",
		X"36",X"01",X"80",X"18",X"12",X"CD",X"39",X"1E",X"30",X"0D",X"CD",X"8E",X"1E",X"DD",X"36",X"00",
		X"00",X"18",X"04",X"FD",X"35",X"01",X"C8",X"3A",X"00",X"4B",X"B7",X"28",X"07",X"3D",X"32",X"00",
		X"4B",X"C3",X"20",X"3C",X"3E",X"00",X"32",X"00",X"4B",X"3A",X"01",X"4B",X"21",X"19",X"3C",X"16",
		X"00",X"5F",X"19",X"7E",X"2A",X"03",X"4B",X"01",X"02",X"05",X"C5",X"E5",X"77",X"23",X"10",X"FC",
		X"E1",X"C1",X"11",X"20",X"00",X"19",X"0D",X"20",X"F1",X"01",X"02",X"05",X"2A",X"05",X"4B",X"C5",
		X"E5",X"77",X"23",X"10",X"FC",X"E1",X"C1",X"11",X"20",X"00",X"19",X"0D",X"20",X"F1",X"2A",X"03",
		X"4B",X"11",X"40",X"00",X"19",X"22",X"03",X"4B",X"2A",X"05",X"4B",X"11",X"C0",X"FF",X"19",X"22",
		X"05",X"4B",X"3A",X"02",X"4B",X"3C",X"FE",X"06",X"38",X"1A",X"11",X"D3",X"45",X"ED",X"53",X"05",
		X"4B",X"21",X"13",X"46",X"22",X"03",X"4B",X"3A",X"01",X"4B",X"3C",X"FE",X"07",X"38",X"01",X"AF",
		X"32",X"01",X"4B",X"AF",X"32",X"02",X"4B",X"18",X"07",X"05",X"04",X"1D",X"17",X"03",X"14",X"15",
		X"3A",X"07",X"4B",X"B7",X"28",X"07",X"3D",X"32",X"07",X"4B",X"C3",X"A1",X"3C",X"3E",X"02",X"32",
		X"07",X"4B",X"3E",X"10",X"CD",X"4B",X"3C",X"3A",X"08",X"4B",X"3C",X"FE",X"04",X"38",X"01",X"AF",
		X"32",X"08",X"4B",X"3E",X"0E",X"CD",X"4B",X"3C",X"C3",X"A1",X"3C",X"F5",X"21",X"78",X"44",X"3A",
		X"08",X"4B",X"06",X"1A",X"B7",X"28",X"07",X"05",X"3D",X"CD",X"79",X"90",X"18",X"F6",X"F1",X"0E",
		X"01",X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"28",X"05",X"CD",X"79",X"90",X"18",X"F2",X"2B",
		X"06",X"06",X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"28",X"03",X"2B",X"18",X"F4",X"11",X"E0",
		X"FF",X"19",X"06",X"19",X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"28",X"06",X"11",X"E0",X"FF",
		X"19",X"18",X"F1",X"23",X"06",X"06",X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"C8",X"23",X"18",
		X"F5",X"3A",X"0A",X"4B",X"FE",X"09",X"D2",X"59",X"3B",X"3A",X"09",X"4B",X"B7",X"28",X"07",X"3D",
		X"32",X"09",X"4B",X"C3",X"59",X"3B",X"3E",X"05",X"32",X"09",X"4B",X"3A",X"0B",X"4B",X"B7",X"20",
		X"16",X"21",X"EB",X"3D",X"CD",X"08",X"3D",X"21",X"3A",X"3E",X"CD",X"08",X"3D",X"3A",X"0B",X"4B",
		X"3C",X"32",X"0B",X"4B",X"C3",X"59",X"3B",X"3A",X"0A",X"4B",X"21",X"EB",X"3D",X"CD",X"1D",X"94",
		X"EB",X"5E",X"23",X"56",X"23",X"EB",X"06",X"1B",X"7E",X"B7",X"28",X"01",X"34",X"CD",X"79",X"90",
		X"10",X"F6",X"3A",X"0B",X"4B",X"3C",X"FE",X"04",X"38",X"08",X"3A",X"0A",X"4B",X"3C",X"32",X"0A",
		X"4B",X"AF",X"32",X"0B",X"4B",X"C3",X"59",X"3B",X"3A",X"0A",X"4B",X"CD",X"1D",X"94",X"EB",X"5E",
		X"23",X"56",X"23",X"EB",X"1A",X"FE",X"FF",X"C8",X"CB",X"7F",X"20",X"0C",X"47",X"13",X"1A",X"77",
		X"CD",X"79",X"90",X"10",X"F8",X"13",X"18",X"EC",X"CB",X"BF",X"47",X"13",X"1A",X"77",X"CD",X"79",
		X"90",X"10",X"FA",X"13",X"C3",X"14",X"3D",X"98",X"40",X"02",X"25",X"5C",X"7E",X"7E",X"7E",X"7F",
		X"80",X"97",X"40",X"02",X"13",X"70",X"71",X"75",X"80",X"B6",X"40",X"02",X"12",X"72",X"76",X"00",
		X"23",X"7E",X"76",X"77",X"80",X"D5",X"40",X"02",X"22",X"73",X"74",X"00",X"31",X"70",X"80",X"38",
		X"41",X"14",X"25",X"5C",X"7E",X"78",X"7E",X"79",X"80",X"37",X"41",X"14",X"13",X"70",X"70",X"75",
		X"00",X"22",X"7E",X"77",X"00",X"32",X"70",X"70",X"80",X"95",X"41",X"14",X"22",X"7C",X"79",X"80",
		X"D8",X"41",X"03",X"25",X"5C",X"7E",X"78",X"7E",X"7F",X"80",X"D7",X"41",X"03",X"13",X"70",X"70",
		X"7D",X"80",X"D5",X"41",X"03",X"12",X"70",X"7D",X"80",X"D3",X"41",X"03",X"13",X"70",X"70",X"7D",
		X"80",X"72",X"42",X"04",X"05",X"79",X"7E",X"78",X"78",X"73",X"00",X"11",X"71",X"00",X"21",X"77",
		X"80",X"B8",X"42",X"04",X"22",X"71",X"72",X"80",X"D8",X"42",X"04",X"25",X"75",X"76",X"76",X"7E",
		X"79",X"80",X"75",X"42",X"04",X"12",X"70",X"70",X"80",X"12",X"43",X"05",X"05",X"79",X"7E",X"7E",
		X"78",X"73",X"00",X"11",X"75",X"00",X"22",X"7A",X"72",X"80",X"54",X"43",X"05",X"03",X"77",X"7A",
		X"73",X"00",X"11",X"75",X"00",X"24",X"76",X"7E",X"7E",X"79",X"FF",X"FD",X"3D",X"0A",X"3E",X"17",
		X"3E",X"1C",X"3E",X"21",X"3E",X"26",X"3E",X"2B",X"3E",X"30",X"3E",X"35",X"3E",X"47",X"40",X"82",
		X"84",X"01",X"8C",X"94",X"00",X"01",X"15",X"83",X"84",X"FF",X"48",X"40",X"84",X"84",X"01",X"8C",
		X"8F",X"00",X"01",X"15",X"86",X"84",X"FF",X"49",X"40",X"9B",X"84",X"FF",X"4A",X"40",X"9B",X"84",
		X"FF",X"4B",X"40",X"9B",X"84",X"FF",X"4C",X"40",X"9B",X"84",X"FF",X"4D",X"40",X"9B",X"84",X"FF",
		X"4E",X"40",X"9B",X"84",X"FF",X"4F",X"40",X"9B",X"84",X"FF",X"4C",X"3E",X"58",X"3E",X"6A",X"3E",
		X"88",X"3E",X"A7",X"3E",X"C5",X"3E",X"E3",X"3E",X"01",X"3F",X"20",X"3F",X"47",X"44",X"83",X"05",
		X"94",X"00",X"04",X"03",X"05",X"03",X"05",X"FF",X"48",X"44",X"83",X"05",X"01",X"03",X"01",X"05",
		X"8F",X"00",X"83",X"05",X"04",X"03",X"05",X"03",X"05",X"FF",X"49",X"44",X"08",X"05",X"03",X"05",
		X"03",X"05",X"03",X"05",X"03",X"83",X"05",X"02",X"03",X"05",X"83",X"03",X"01",X"05",X"83",X"03",
		X"83",X"05",X"04",X"03",X"05",X"03",X"05",X"FF",X"4A",X"44",X"0D",X"03",X"03",X"05",X"03",X"05",
		X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"83",X"03",X"01",X"05",X"83",X"03",X"01",X"05",
		X"83",X"03",X"03",X"05",X"03",X"05",X"FF",X"4B",X"44",X"83",X"05",X"0A",X"03",X"05",X"03",X"05",
		X"03",X"05",X"03",X"05",X"03",X"05",X"83",X"03",X"01",X"05",X"83",X"03",X"01",X"05",X"83",X"03",
		X"03",X"05",X"05",X"03",X"FF",X"4C",X"44",X"01",X"05",X"83",X"03",X"83",X"05",X"05",X"03",X"05",
		X"03",X"05",X"03",X"83",X"05",X"01",X"03",X"83",X"05",X"01",X"03",X"83",X"05",X"04",X"03",X"05",
		X"03",X"05",X"FF",X"4D",X"44",X"01",X"05",X"83",X"03",X"83",X"05",X"0E",X"03",X"05",X"03",X"05",
		X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"83",X"03",X"03",X"05",X"03",X"05",
		X"FF",X"4E",X"44",X"15",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",
		X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"03",X"05",X"83",X"03",X"03",X"05",X"03",X"05",X"FF",
		X"4F",X"44",X"83",X"05",X"05",X"03",X"05",X"03",X"05",X"03",X"83",X"05",X"01",X"03",X"83",X"05",
		X"01",X"03",X"83",X"05",X"01",X"03",X"83",X"05",X"01",X"03",X"83",X"05",X"FF",X"FF",X"FF",X"FF",
		X"31",X"E0",X"4D",X"21",X"C0",X"4A",X"06",X"0F",X"CF",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",
		X"C0",X"4A",X"06",X"05",X"C5",X"FD",X"7E",X"00",X"B7",X"28",X"06",X"FD",X"35",X"00",X"CC",X"6B",
		X"3F",X"01",X"03",X"00",X"FD",X"09",X"C1",X"10",X"EB",X"18",X"DE",X"FD",X"7E",X"01",X"CD",X"EA",
		X"91",X"CD",X"1E",X"92",X"CD",X"83",X"26",X"38",X"10",X"E5",X"FD",X"7E",X"02",X"E6",X"07",X"CD",
		X"87",X"95",X"E1",X"01",X"02",X"02",X"CD",X"5C",X"90",X"FD",X"E5",X"E1",X"06",X"03",X"CF",X"C9",
		X"FD",X"E5",X"FD",X"21",X"C0",X"4A",X"06",X"05",X"FD",X"7E",X"00",X"B7",X"28",X"0D",X"FD",X"23",
		X"FD",X"23",X"FD",X"23",X"10",X"F2",X"FD",X"E1",X"C9",X"10",X"ED",X"01",X"68",X"48",X"7E",X"B7",
		X"ED",X"42",X"FD",X"36",X"00",X"12",X"FD",X"75",X"01",X"FD",X"77",X"02",X"FD",X"E1",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
