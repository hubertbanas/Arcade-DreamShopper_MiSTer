library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"E0",X"4E",X"3A",X"AA",X"49",X"FE",X"03",X"30",X"03",X"3E",X"60",X"FF",X"21",X"45",X"48",
		X"06",X"0A",X"CF",X"21",X"00",X"4A",X"06",X"20",X"CF",X"FD",X"21",X"00",X"4A",X"CD",X"A6",X"82",
		X"FD",X"21",X"10",X"4A",X"CD",X"A6",X"82",X"29",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"3E",X"23",
		X"06",X"01",X"FF",X"FD",X"21",X"00",X"4A",X"DD",X"21",X"45",X"48",X"CD",X"AB",X"85",X"3A",X"01",
		X"48",X"CB",X"47",X"28",X"2E",X"DD",X"E5",X"E1",X"06",X"0A",X"CF",X"3E",X"23",X"06",X"01",X"FF",
		X"3A",X"01",X"48",X"CB",X"47",X"20",X"F4",X"11",X"46",X"48",X"21",X"03",X"4A",X"01",X"04",X"00",
		X"ED",X"B0",X"11",X"4B",X"48",X"21",X"13",X"4A",X"01",X"04",X"00",X"ED",X"B0",X"DD",X"36",X"00",
		X"01",X"18",X"BB",X"C5",X"FD",X"7E",X"00",X"E6",X"0F",X"21",X"8C",X"80",X"E5",X"DF",X"B1",X"80",
		X"CB",X"81",X"34",X"81",X"45",X"81",X"56",X"81",X"94",X"81",X"64",X"81",X"DD",X"E5",X"E1",X"23",
		X"FD",X"E5",X"D1",X"13",X"13",X"13",X"01",X"04",X"00",X"ED",X"B0",X"DD",X"36",X"00",X"00",X"01",
		X"05",X"00",X"DD",X"09",X"01",X"10",X"00",X"FD",X"09",X"C1",X"05",X"C2",X"73",X"80",X"C3",X"2E",
		X"80",X"FD",X"6E",X"0E",X"FD",X"66",X"0F",X"7D",X"B4",X"28",X"08",X"2B",X"FD",X"75",X"0E",X"FD",
		X"74",X"0F",X"C9",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"05",X"3E",X"15",X"C3",X"03",X"81",X"11",
		X"00",X"00",X"21",X"68",X"48",X"ED",X"5F",X"E6",X"7F",X"06",X"00",X"4F",X"09",X"7E",X"FE",X"03",
		X"28",X"18",X"23",X"E5",X"01",X"F8",X"48",X"AF",X"ED",X"42",X"E1",X"20",X"F0",X"3C",X"BA",X"28",
		X"06",X"14",X"21",X"68",X"48",X"18",X"E6",X"3E",X"60",X"FF",X"CB",X"DE",X"AF",X"01",X"68",X"48",
		X"ED",X"42",X"7D",X"CD",X"EA",X"91",X"DD",X"36",X"01",X"18",X"DD",X"74",X"02",X"DD",X"36",X"03",
		X"16",X"DD",X"75",X"04",X"DD",X"36",X"00",X"00",X"CD",X"1E",X"92",X"3E",X"29",X"1E",X"51",X"01",
		X"02",X"02",X"CD",X"5C",X"90",X"FD",X"36",X"00",X"01",X"FD",X"36",X"07",X"0A",X"CD",X"A6",X"82",
		X"CD",X"83",X"82",X"C9",X"FD",X"CB",X"00",X"76",X"C2",X"88",X"85",X"FD",X"7E",X"08",X"B7",X"C2",
		X"46",X"82",X"C3",X"72",X"84",X"FD",X"CB",X"00",X"76",X"C2",X"88",X"85",X"FD",X"7E",X"08",X"B7",
		X"C2",X"46",X"82",X"C3",X"CE",X"82",X"FD",X"CB",X"00",X"6E",X"28",X"03",X"C3",X"9E",X"85",X"CD",
		X"7A",X"81",X"18",X"E1",X"FD",X"CB",X"00",X"6E",X"28",X"03",X"C3",X"9E",X"85",X"CD",X"7A",X"81",
		X"FD",X"7E",X"08",X"B7",X"C2",X"46",X"82",X"C3",X"94",X"83",X"FD",X"7E",X"07",X"B7",X"20",X"10",
		X"FD",X"36",X"07",X"06",X"3E",X"36",X"DD",X"BE",X"01",X"20",X"02",X"3E",X"37",X"DD",X"77",X"01",
		X"FD",X"35",X"07",X"C9",X"FD",X"7E",X"07",X"B7",X"28",X"02",X"18",X"10",X"FD",X"36",X"07",X"06",
		X"3E",X"37",X"DD",X"BE",X"01",X"20",X"02",X"3E",X"38",X"DD",X"77",X"01",X"FD",X"35",X"07",X"FD",
		X"7E",X"08",X"B7",X"C2",X"46",X"82",X"21",X"00",X"02",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",
		X"FF",X"FF",X"FD",X"75",X"01",X"FD",X"74",X"02",X"C3",X"46",X"82",X"FD",X"7E",X"07",X"B7",X"28",
		X"04",X"FD",X"35",X"07",X"C9",X"DD",X"34",X"01",X"3E",X"1E",X"DD",X"BE",X"01",X"28",X"05",X"FD",
		X"36",X"07",X"0A",X"C9",X"DD",X"36",X"01",X"36",X"DD",X"36",X"03",X"51",X"DD",X"66",X"02",X"DD",
		X"6E",X"04",X"E5",X"CD",X"AC",X"91",X"CB",X"9E",X"CB",X"7E",X"E1",X"20",X"0D",X"CD",X"1E",X"92",
		X"01",X"02",X"02",X"1E",X"16",X"3E",X"00",X"CD",X"0C",X"90",X"DD",X"7E",X"04",X"FD",X"36",X"00",
		X"03",X"FE",X"50",X"38",X"04",X"FD",X"36",X"00",X"02",X"FD",X"CB",X"00",X"FE",X"DD",X"7E",X"02",
		X"FE",X"88",X"D0",X"FD",X"CB",X"00",X"BE",X"C9",X"FD",X"6E",X"01",X"FD",X"66",X"02",X"29",X"38",
		X"07",X"FD",X"75",X"01",X"FD",X"74",X"02",X"C9",X"F5",X"11",X"00",X"00",X"ED",X"5A",X"FD",X"75",
		X"01",X"FD",X"74",X"02",X"F1",X"C9",X"CD",X"28",X"82",X"D0",X"FD",X"4E",X"09",X"FD",X"46",X"0A",
		X"DD",X"66",X"02",X"DD",X"6E",X"04",X"FD",X"CB",X"00",X"7E",X"28",X"04",X"79",X"ED",X"44",X"4F",
		X"CD",X"A5",X"91",X"DD",X"74",X"02",X"DD",X"75",X"04",X"FD",X"35",X"08",X"DD",X"7E",X"04",X"FE",
		X"02",X"C0",X"DD",X"E5",X"E1",X"06",X"05",X"CF",X"FD",X"E5",X"E1",X"06",X"0E",X"CF",X"DD",X"36",
		X"00",X"00",X"C9",X"21",X"9A",X"82",X"3A",X"AA",X"49",X"FE",X"06",X"38",X"02",X"3E",X"06",X"3D",
		X"CD",X"1D",X"94",X"FD",X"73",X"01",X"FD",X"72",X"02",X"C9",X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",
		X"D6",X"D6",X"AA",X"AA",X"EE",X"EE",X"3A",X"AA",X"49",X"FE",X"08",X"38",X"02",X"3E",X"08",X"3D",
		X"21",X"BE",X"82",X"CD",X"1D",X"94",X"EB",X"FD",X"75",X"0E",X"FD",X"74",X"0F",X"C9",X"5A",X"02",
		X"5A",X"02",X"E1",X"01",X"70",X"01",X"30",X"01",X"F0",X"00",X"B4",X"00",X"78",X"00",X"FD",X"6E",
		X"0B",X"FD",X"66",X"0C",X"7D",X"B4",X"28",X"2B",X"7E",X"FE",X"FF",X"28",X"15",X"23",X"5E",X"23",
		X"56",X"23",X"FD",X"77",X"09",X"FD",X"73",X"0A",X"FD",X"72",X"08",X"FD",X"75",X"0B",X"FD",X"74",
		X"0C",X"C9",X"3A",X"2C",X"48",X"CB",X"7F",X"20",X"0A",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"06",
		X"CD",X"40",X"03",X"FD",X"7E",X"00",X"E6",X"0F",X"FE",X"04",X"C2",X"3C",X"85",X"06",X"03",X"3A",
		X"AA",X"49",X"FE",X"05",X"38",X"02",X"06",X"00",X"FD",X"7E",X"0D",X"B8",X"DA",X"B7",X"83",X"3A",
		X"42",X"48",X"C6",X"F0",X"5F",X"C6",X"20",X"57",X"DD",X"7E",X"02",X"BB",X"DA",X"B7",X"83",X"BA",
		X"D2",X"B7",X"83",X"DD",X"7E",X"02",X"E6",X"0F",X"CA",X"94",X"83",X"FD",X"36",X"00",X"06",X"DD",
		X"5E",X"02",X"3A",X"42",X"48",X"93",X"28",X"1C",X"30",X"0B",X"DD",X"7E",X"02",X"E6",X"0F",X"FD",
		X"CB",X"00",X"FE",X"18",X"1A",X"DD",X"7E",X"02",X"E6",X"0F",X"ED",X"44",X"E6",X"0F",X"FD",X"CB",
		X"00",X"BE",X"18",X"0B",X"DD",X"7E",X"02",X"E6",X"0F",X"CB",X"5F",X"28",X"DD",X"18",X"E6",X"FD",
		X"CB",X"00",X"EE",X"FD",X"77",X"08",X"FD",X"36",X"07",X"04",X"DD",X"36",X"01",X"36",X"21",X"01",
		X"00",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"00",X"00",X"FD",X"75",X"0B",X"FD",X"74",X"0C",
		X"CD",X"83",X"82",X"C9",X"21",X"00",X"FF",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"FD",X"36",X"08",
		X"00",X"DD",X"36",X"01",X"37",X"FD",X"36",X"00",X"05",X"FD",X"36",X"07",X"06",X"CD",X"9A",X"2D",
		X"C8",X"3E",X"07",X"CD",X"40",X"03",X"C9",X"06",X"05",X"3E",X"48",X"0E",X"00",X"DD",X"BE",X"04",
		X"30",X"0C",X"C6",X"10",X"F5",X"79",X"C6",X"08",X"4F",X"F1",X"10",X"F1",X"0E",X"20",X"06",X"00",
		X"21",X"25",X"08",X"09",X"ED",X"5F",X"E6",X"03",X"CD",X"1D",X"94",X"EB",X"06",X"00",X"7E",X"FD",
		X"CB",X"00",X"7E",X"28",X"22",X"ED",X"44",X"5F",X"16",X"FF",X"E5",X"DD",X"6E",X"02",X"26",X"00",
		X"19",X"7D",X"E1",X"30",X"04",X"FE",X"30",X"30",X"30",X"3E",X"01",X"B8",X"CA",X"30",X"85",X"06",
		X"01",X"FD",X"CB",X"00",X"BE",X"18",X"D7",X"E5",X"DD",X"6E",X"02",X"26",X"00",X"5F",X"16",X"00",
		X"19",X"7D",X"CB",X"44",X"E1",X"20",X"04",X"FE",X"E1",X"38",X"0E",X"3E",X"01",X"B8",X"CA",X"30",
		X"85",X"06",X"01",X"FD",X"CB",X"00",X"FE",X"18",X"B5",X"FD",X"7E",X"00",X"E6",X"80",X"F6",X"03",
		X"FD",X"77",X"00",X"FD",X"34",X"0D",X"23",X"4E",X"23",X"46",X"23",X"56",X"23",X"5E",X"23",X"7E",
		X"23",X"FD",X"75",X"0B",X"FD",X"74",X"0C",X"FD",X"72",X"09",X"FD",X"73",X"0A",X"FD",X"77",X"08",
		X"FD",X"71",X"01",X"FD",X"70",X"02",X"FD",X"36",X"07",X"04",X"FD",X"CB",X"00",X"F6",X"DD",X"36",
		X"01",X"36",X"3A",X"2C",X"48",X"CB",X"7F",X"C0",X"CD",X"9A",X"2D",X"C8",X"3E",X"06",X"CD",X"40",
		X"03",X"C9",X"FD",X"6E",X"0B",X"FD",X"66",X"0C",X"7D",X"B4",X"28",X"3A",X"7E",X"FE",X"FF",X"28",
		X"15",X"23",X"5E",X"23",X"56",X"23",X"FD",X"77",X"09",X"FD",X"73",X"0A",X"FD",X"72",X"08",X"FD",
		X"75",X"0B",X"FD",X"74",X"0C",X"C9",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"06",X"CD",X"40",X"03",
		X"21",X"00",X"00",X"FD",X"75",X"0B",X"FD",X"74",X"0C",X"FD",X"CB",X"00",X"EE",X"FD",X"36",X"07",
		X"04",X"DD",X"36",X"01",X"36",X"C9",X"21",X"AB",X"09",X"ED",X"5F",X"E6",X"03",X"CD",X"17",X"94",
		X"5E",X"23",X"56",X"EB",X"7E",X"23",X"DD",X"86",X"04",X"FE",X"40",X"30",X"12",X"21",X"00",X"00",
		X"FD",X"75",X"0B",X"FD",X"74",X"0C",X"FD",X"36",X"08",X"00",X"FD",X"36",X"00",X"03",X"C9",X"06",
		X"00",X"7E",X"FD",X"CB",X"00",X"7E",X"28",X"26",X"ED",X"44",X"5F",X"16",X"FF",X"E5",X"DD",X"6E",
		X"02",X"26",X"00",X"19",X"7D",X"E1",X"30",X"09",X"DD",X"7E",X"02",X"83",X"FE",X"30",X"D2",X"36",
		X"84",X"3E",X"01",X"B8",X"28",X"2A",X"06",X"01",X"FD",X"CB",X"00",X"BE",X"18",X"D3",X"E5",X"DD",
		X"6E",X"02",X"26",X"00",X"16",X"00",X"5F",X"19",X"7D",X"CB",X"44",X"E1",X"20",X"05",X"FE",X"E1",
		X"DA",X"36",X"84",X"3E",X"01",X"B8",X"28",X"08",X"06",X"01",X"FD",X"CB",X"00",X"FE",X"18",X"B1",
		X"21",X"36",X"85",X"C3",X"37",X"84",X"AA",X"AA",X"00",X"00",X"08",X"FF",X"ED",X"5F",X"E6",X"1F",
		X"C6",X"10",X"5F",X"DD",X"7E",X"02",X"FD",X"CB",X"00",X"7E",X"FD",X"36",X"00",X"04",X"28",X"2B",
		X"93",X"FE",X"30",X"38",X"2D",X"FD",X"CB",X"00",X"FE",X"DD",X"36",X"01",X"36",X"FD",X"73",X"08",
		X"21",X"01",X"00",X"FD",X"75",X"09",X"FD",X"74",X"0A",X"21",X"00",X"00",X"FD",X"75",X"0B",X"FD",
		X"74",X"0C",X"FD",X"CB",X"00",X"EE",X"FD",X"36",X"07",X"04",X"C9",X"83",X"38",X"D7",X"FE",X"E1",
		X"30",X"D3",X"DD",X"36",X"01",X"36",X"18",X"D5",X"FD",X"35",X"07",X"C0",X"3E",X"9F",X"FD",X"A6",
		X"00",X"FD",X"CB",X"00",X"76",X"FD",X"77",X"00",X"C8",X"DD",X"36",X"01",X"38",X"C9",X"FD",X"35",
		X"07",X"C0",X"FD",X"CB",X"00",X"AE",X"DD",X"36",X"01",X"36",X"C9",X"3A",X"AA",X"49",X"FE",X"06",
		X"38",X"02",X"3E",X"06",X"3D",X"21",X"BE",X"85",X"16",X"00",X"5F",X"19",X"46",X"C9",X"01",X"01",
		X"01",X"01",X"01",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"20",X"4F",X"21",X"4A",X"48",X"06",X"14",X"CF",X"21",X"20",X"4A",X"06",X"3F",X"CF",X"CD",
		X"70",X"89",X"0E",X"00",X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"04",X"D6",X"09",X"18",X"F8",X"FE",
		X"04",X"38",X"05",X"D6",X"03",X"0C",X"18",X"F7",X"3D",X"32",X"24",X"4A",X"79",X"32",X"23",X"4A",
		X"3E",X"23",X"06",X"01",X"FF",X"CD",X"C4",X"8A",X"FD",X"21",X"27",X"4A",X"DD",X"21",X"4F",X"48",
		X"CD",X"91",X"8E",X"21",X"97",X"49",X"3A",X"01",X"48",X"CB",X"47",X"28",X"30",X"DD",X"E5",X"E1",
		X"06",X"14",X"CF",X"3E",X"23",X"06",X"01",X"FF",X"3A",X"01",X"48",X"CB",X"47",X"20",X"F4",X"11",
		X"04",X"00",X"FD",X"19",X"11",X"4F",X"48",X"06",X"04",X"C5",X"FD",X"E5",X"E1",X"13",X"01",X"04",
		X"00",X"ED",X"B0",X"01",X"0E",X"00",X"FD",X"09",X"C1",X"10",X"EE",X"18",X"B3",X"C5",X"E5",X"FD",
		X"7E",X"00",X"E6",X"0F",X"B7",X"CA",X"57",X"87",X"3D",X"21",X"96",X"86",X"E5",X"DF",X"BB",X"87",
		X"FD",X"87",X"FD",X"87",X"CC",X"88",X"FD",X"7E",X"00",X"B7",X"28",X"15",X"FE",X"04",X"30",X"11",
		X"FD",X"7E",X"08",X"B7",X"28",X"05",X"FD",X"35",X"08",X"18",X"06",X"CD",X"29",X"89",X"CD",X"E6",
		X"8B",X"DD",X"E5",X"D1",X"13",X"FD",X"E5",X"E1",X"23",X"23",X"23",X"23",X"01",X"04",X"00",X"ED",
		X"B0",X"DD",X"36",X"00",X"00",X"E1",X"23",X"23",X"11",X"05",X"00",X"DD",X"19",X"11",X"0E",X"00",
		X"FD",X"19",X"C1",X"05",X"C2",X"7D",X"86",X"3A",X"20",X"4A",X"B7",X"20",X"11",X"ED",X"5F",X"32",
		X"20",X"4A",X"F5",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"11",X"CD",X"40",X"03",X"F1",X"3D",X"32",
		X"20",X"4A",X"2A",X"25",X"4A",X"7D",X"B4",X"CA",X"30",X"86",X"2B",X"7D",X"B4",X"28",X"33",X"AF",
		X"B4",X"20",X"29",X"7D",X"FE",X"40",X"30",X"24",X"E6",X"03",X"20",X"20",X"FD",X"21",X"27",X"4A",
		X"06",X"05",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"0C",X"3E",X"53",X"FD",X"BE",X"06",X"20",X"02",
		X"3E",X"52",X"FD",X"77",X"06",X"11",X"0E",X"00",X"FD",X"19",X"10",X"E6",X"22",X"25",X"4A",X"C3",
		X"30",X"86",X"FD",X"21",X"27",X"4A",X"06",X"05",X"FD",X"7E",X"00",X"FE",X"02",X"20",X"0E",X"C5",
		X"3E",X"84",X"CD",X"40",X"03",X"C1",X"FD",X"36",X"00",X"03",X"CD",X"03",X"89",X"11",X"0E",X"00",
		X"FD",X"19",X"10",X"E4",X"C3",X"30",X"86",X"5E",X"23",X"56",X"7B",X"B2",X"28",X"07",X"1B",X"72",
		X"2B",X"73",X"C3",X"96",X"86",X"11",X"00",X"01",X"72",X"2B",X"73",X"21",X"F9",X"8D",X"3A",X"21",
		X"4A",X"E6",X"03",X"CD",X"16",X"94",X"7E",X"23",X"56",X"23",X"5E",X"23",X"4E",X"FD",X"77",X"01",
		X"FD",X"71",X"09",X"FD",X"72",X"05",X"FD",X"73",X"07",X"CD",X"03",X"89",X"CD",X"09",X"8E",X"CD",
		X"4D",X"8E",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"16",X"3A",X"21",X"4A",X"21",X"4D",X"0A",X"CD",
		X"17",X"94",X"5E",X"23",X"56",X"FD",X"73",X"0A",X"FD",X"72",X"0B",X"3E",X"03",X"18",X"02",X"3E",
		X"01",X"FD",X"77",X"00",X"21",X"21",X"4A",X"34",X"C3",X"96",X"86",X"FD",X"5E",X"0A",X"FD",X"56",
		X"0B",X"7B",X"B2",X"28",X"07",X"1B",X"FD",X"73",X"0A",X"FD",X"72",X"0B",X"CD",X"19",X"8B",X"D0",
		X"CD",X"37",X"8B",X"C2",X"DD",X"88",X"CD",X"6D",X"8D",X"5F",X"FD",X"7E",X"01",X"E6",X"03",X"CD",
		X"31",X"94",X"A3",X"CA",X"04",X"8C",X"FD",X"7E",X"09",X"B7",X"C2",X"DD",X"88",X"FD",X"5E",X"0A",
		X"FD",X"56",X"0B",X"7B",X"B2",X"C2",X"04",X"8C",X"FD",X"36",X"00",X"03",X"C9",X"3A",X"02",X"48",
		X"CB",X"77",X"28",X"75",X"FD",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"FD",X"21",X"A0",X"4A",
		X"06",X"03",X"FD",X"7E",X"00",X"FE",X"02",X"C2",X"6E",X"88",X"FD",X"7E",X"03",X"C6",X"F8",X"57",
		X"C6",X"50",X"5F",X"DD",X"7E",X"05",X"BA",X"DA",X"6E",X"88",X"BB",X"D2",X"6E",X"88",X"FD",X"7E",
		X"04",X"C6",X"B8",X"57",X"C6",X"50",X"5F",X"DD",X"7E",X"07",X"BA",X"38",X"31",X"BB",X"30",X"2E",
		X"DD",X"E1",X"FD",X"E1",X"CD",X"9A",X"2D",X"28",X"05",X"3E",X"0C",X"CD",X"40",X"03",X"FD",X"36",
		X"00",X"04",X"FD",X"36",X"01",X"40",X"FD",X"36",X"06",X"03",X"FD",X"36",X"04",X"35",X"21",X"6D",
		X"88",X"CD",X"BA",X"2C",X"C2",X"D5",X"2C",X"C9",X"00",X"00",X"00",X"01",X"00",X"00",X"11",X"0A",
		X"00",X"FD",X"19",X"10",X"9D",X"DD",X"E1",X"FD",X"E1",X"CD",X"19",X"8B",X"D0",X"3E",X"03",X"FD",
		X"BE",X"00",X"20",X"07",X"FD",X"CB",X"01",X"6E",X"C4",X"F6",X"8C",X"CD",X"37",X"8B",X"C2",X"DD",
		X"88",X"3A",X"01",X"48",X"CB",X"7F",X"CA",X"9C",X"8E",X"FD",X"7E",X"00",X"E6",X"0F",X"FE",X"02",
		X"1E",X"0F",X"20",X"04",X"CD",X"C4",X"8E",X"5F",X"D5",X"CD",X"B5",X"8D",X"D1",X"A3",X"5F",X"D5",
		X"CD",X"94",X"8D",X"D1",X"A3",X"5F",X"FD",X"7E",X"01",X"E6",X"03",X"CD",X"31",X"94",X"A3",X"CA",
		X"2C",X"8C",X"FD",X"7E",X"09",X"B7",X"CA",X"2C",X"8C",X"C3",X"DD",X"88",X"FD",X"35",X"01",X"C0",
		X"DD",X"E5",X"E1",X"06",X"05",X"CF",X"FD",X"E5",X"E1",X"06",X"0E",X"CF",X"C9",X"FD",X"35",X"09",
		X"21",X"89",X"8E",X"FD",X"7E",X"01",X"E6",X"03",X"CD",X"17",X"94",X"4E",X"23",X"46",X"FD",X"66",
		X"05",X"FD",X"6E",X"07",X"CD",X"A5",X"91",X"FD",X"74",X"05",X"FD",X"75",X"07",X"C9",X"21",X"19",
		X"89",X"18",X"03",X"21",X"21",X"89",X"FD",X"7E",X"01",X"E6",X"03",X"CD",X"1D",X"94",X"FD",X"73",
		X"04",X"FD",X"72",X"06",X"FD",X"CB",X"01",X"BE",X"C9",X"30",X"53",X"AD",X"53",X"30",X"53",X"2D",
		X"53",X"2B",X"52",X"A8",X"52",X"2B",X"52",X"28",X"52",X"21",X"68",X"89",X"3E",X"02",X"FD",X"BE",
		X"00",X"28",X"03",X"21",X"60",X"89",X"FD",X"7E",X"01",X"E6",X"03",X"CD",X"1D",X"94",X"FD",X"CB",
		X"01",X"7E",X"20",X"0E",X"7A",X"FD",X"BE",X"04",X"28",X"0E",X"FD",X"CB",X"01",X"BE",X"FD",X"34",
		X"04",X"C9",X"7B",X"FD",X"BE",X"04",X"28",X"F2",X"FD",X"CB",X"01",X"FE",X"FD",X"35",X"04",X"C9",
		X"2B",X"2C",X"A8",X"AA",X"2B",X"2C",X"28",X"2A",X"30",X"31",X"AD",X"AF",X"30",X"31",X"2D",X"2F",
		X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"5F",X"87",X"83",X"5F",X"3A",X"A4",
		X"49",X"FE",X"02",X"38",X"02",X"3E",X"02",X"83",X"21",X"98",X"89",X"CD",X"1D",X"94",X"EB",X"11",
		X"97",X"49",X"01",X"08",X"00",X"ED",X"B0",X"C9",X"D4",X"89",X"DC",X"89",X"E4",X"89",X"EC",X"89",
		X"F4",X"89",X"FC",X"89",X"04",X"8A",X"0C",X"8A",X"14",X"8A",X"1C",X"8A",X"24",X"8A",X"2C",X"8A",
		X"34",X"8A",X"3C",X"8A",X"44",X"8A",X"4C",X"8A",X"54",X"8A",X"5C",X"8A",X"64",X"8A",X"6C",X"8A",
		X"74",X"8A",X"7C",X"8A",X"84",X"8A",X"8C",X"8A",X"94",X"8A",X"9C",X"8A",X"A4",X"8A",X"AC",X"8A",
		X"B4",X"8A",X"BC",X"8A",X"F0",X"00",X"58",X"02",X"84",X"03",X"B0",X"04",X"00",X"00",X"2C",X"01",
		X"58",X"02",X"84",X"03",X"00",X"00",X"00",X"00",X"58",X"02",X"84",X"03",X"B4",X"00",X"E0",X"01",
		X"D0",X"02",X"84",X"03",X"00",X"00",X"F0",X"00",X"E0",X"01",X"D0",X"02",X"00",X"00",X"00",X"00",
		X"E0",X"01",X"D0",X"02",X"B4",X"00",X"2C",X"01",X"58",X"02",X"84",X"03",X"00",X"00",X"F0",X"00",
		X"F0",X"00",X"58",X"02",X"00",X"00",X"00",X"00",X"F0",X"00",X"58",X"02",X"F0",X"00",X"E0",X"01",
		X"D0",X"02",X"84",X"03",X"00",X"00",X"F0",X"00",X"E0",X"01",X"D0",X"02",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"E0",X"01",X"B4",X"00",X"68",X"01",X"D0",X"02",X"D0",X"02",X"00",X"00",X"68",X"01",
		X"D0",X"02",X"84",X"03",X"00",X"00",X"00",X"00",X"68",X"01",X"D0",X"02",X"B4",X"00",X"84",X"03",
		X"D0",X"05",X"08",X"07",X"00",X"00",X"2C",X"01",X"58",X"02",X"84",X"03",X"00",X"00",X"00",X"00",
		X"2C",X"01",X"58",X"02",X"B4",X"00",X"E0",X"01",X"D0",X"02",X"B0",X"04",X"00",X"00",X"B4",X"00",
		X"E0",X"01",X"58",X"02",X"00",X"00",X"00",X"00",X"B4",X"00",X"E0",X"01",X"B4",X"00",X"2C",X"01",
		X"2C",X"01",X"2C",X"01",X"00",X"00",X"2C",X"01",X"58",X"02",X"84",X"03",X"00",X"00",X"00",X"00",
		X"2C",X"01",X"58",X"02",X"B4",X"00",X"B4",X"00",X"2C",X"01",X"58",X"02",X"00",X"00",X"B4",X"00",
		X"2C",X"01",X"58",X"02",X"00",X"00",X"00",X"00",X"B4",X"00",X"2C",X"01",X"00",X"00",X"00",X"00",
		X"58",X"02",X"84",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"58",X"02",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"21",X"F6",X"8A",X"3A",X"AA",X"49",X"FE",X"02",X"30",X"03",X"21",X"FC",
		X"8A",X"0E",X"00",X"E5",X"06",X"02",X"11",X"94",X"49",X"CD",X"80",X"90",X"E1",X"FE",X"01",X"28",
		X"0E",X"0C",X"79",X"FE",X"03",X"38",X"04",X"0E",X"02",X"18",X"04",X"23",X"23",X"18",X"E4",X"79",
		X"21",X"24",X"4A",X"86",X"77",X"C9",X"1E",X"00",X"28",X"00",X"3C",X"00",X"1E",X"00",X"3C",X"00",
		X"3C",X"00",X"3A",X"24",X"4A",X"FE",X"04",X"38",X"02",X"3E",X"04",X"21",X"14",X"8B",X"16",X"00",
		X"5F",X"19",X"7E",X"C9",X"20",X"10",X"08",X"08",X"08",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"29",
		X"38",X"07",X"FD",X"75",X"02",X"FD",X"74",X"03",X"C9",X"F5",X"11",X"00",X"00",X"ED",X"5A",X"FD",
		X"75",X"02",X"FD",X"74",X"03",X"F1",X"C9",X"FD",X"7E",X"05",X"E6",X"0F",X"C0",X"FD",X"7E",X"07",
		X"E6",X"0F",X"C0",X"C9",X"CD",X"24",X"94",X"21",X"86",X"8B",X"F5",X"FD",X"7E",X"00",X"FE",X"02",
		X"28",X"03",X"21",X"B6",X"8B",X"F1",X"CD",X"16",X"94",X"FD",X"7E",X"01",X"E6",X"70",X"B6",X"FD",
		X"77",X"01",X"23",X"7E",X"FD",X"77",X"04",X"3A",X"01",X"48",X"CB",X"7F",X"28",X"14",X"23",X"5E",
		X"23",X"56",X"EB",X"ED",X"5F",X"E6",X"07",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",X"09",X"CD",
		X"DD",X"88",X"CD",X"E6",X"8B",X"C9",X"00",X"30",X"96",X"8B",X"01",X"AD",X"9E",X"8B",X"02",X"30",
		X"A6",X"8B",X"03",X"2D",X"AE",X"8B",X"40",X"20",X"50",X"40",X"10",X"30",X"40",X"20",X"30",X"50",
		X"40",X"20",X"10",X"40",X"30",X"20",X"40",X"20",X"30",X"40",X"50",X"10",X"40",X"30",X"30",X"50",
		X"20",X"40",X"10",X"40",X"30",X"20",X"00",X"2B",X"C6",X"8B",X"01",X"A8",X"CE",X"8B",X"02",X"2B",
		X"D6",X"8B",X"03",X"28",X"DE",X"8B",X"30",X"20",X"50",X"10",X"20",X"10",X"10",X"30",X"10",X"30",
		X"40",X"20",X"10",X"30",X"20",X"10",X"30",X"20",X"10",X"40",X"50",X"10",X"20",X"10",X"20",X"10",
		X"30",X"40",X"10",X"40",X"30",X"10",X"21",X"FC",X"8B",X"3A",X"AA",X"49",X"3D",X"FE",X"07",X"38",
		X"02",X"3E",X"07",X"16",X"00",X"5F",X"19",X"7E",X"FD",X"77",X"08",X"C9",X"05",X"04",X"03",X"03",
		X"03",X"03",X"03",X"03",X"CD",X"B5",X"8D",X"1E",X"0F",X"A3",X"5F",X"D5",X"CD",X"6D",X"8D",X"D1",
		X"A3",X"5F",X"ED",X"5F",X"E6",X"03",X"CD",X"31",X"94",X"A3",X"C8",X"4F",X"3A",X"96",X"49",X"FE",
		X"02",X"79",X"DA",X"44",X"8B",X"3E",X"0E",X"A3",X"C8",X"C3",X"44",X"8B",X"FD",X"7E",X"00",X"E6",
		X"0F",X"FE",X"02",X"CA",X"23",X"8D",X"3A",X"E9",X"49",X"E6",X"07",X"FE",X"04",X"38",X"0E",X"FD",
		X"CB",X"01",X"76",X"FD",X"CB",X"01",X"F6",X"28",X"68",X"FD",X"CB",X"01",X"B6",X"FD",X"CB",X"01",
		X"46",X"28",X"13",X"1E",X"04",X"3A",X"44",X"48",X"B7",X"28",X"19",X"FD",X"BE",X"07",X"28",X"06",
		X"30",X"12",X"1E",X"01",X"18",X"0E",X"1E",X"02",X"3A",X"42",X"48",X"FD",X"BE",X"05",X"28",X"E3",
		X"30",X"02",X"1E",X"08",X"3A",X"44",X"48",X"FD",X"BE",X"07",X"28",X"13",X"3A",X"42",X"48",X"FD",
		X"BE",X"05",X"28",X"0B",X"FD",X"CB",X"01",X"AE",X"D5",X"CD",X"09",X"8E",X"D1",X"18",X"12",X"FD",
		X"CB",X"01",X"EE",X"20",X"0C",X"FD",X"36",X"0C",X"00",X"D5",X"CD",X"02",X"8B",X"FD",X"77",X"0D",
		X"D1",X"D5",X"CD",X"B5",X"8D",X"D1",X"A3",X"5F",X"D5",X"CD",X"94",X"8D",X"D1",X"A3",X"C2",X"44",
		X"8B",X"1E",X"0F",X"D5",X"CD",X"B5",X"8D",X"D1",X"A3",X"5F",X"D5",X"CD",X"94",X"8D",X"D1",X"A3",
		X"CA",X"04",X"8C",X"5F",X"ED",X"5F",X"E6",X"07",X"47",X"ED",X"5F",X"CB",X"07",X"10",X"FC",X"E6",
		X"03",X"CD",X"31",X"94",X"A3",X"C8",X"5F",X"3E",X"05",X"FD",X"CB",X"01",X"46",X"20",X"02",X"3E",
		X"0A",X"A3",X"C2",X"44",X"8B",X"FD",X"CB",X"01",X"66",X"FD",X"CB",X"01",X"E6",X"C8",X"FD",X"CB",
		X"01",X"A6",X"7B",X"C3",X"44",X"8B",X"FD",X"7E",X"0D",X"B7",X"28",X"04",X"FD",X"35",X"0D",X"C9",
		X"FD",X"7E",X"0C",X"FE",X"03",X"C8",X"FD",X"36",X"0D",X"08",X"3C",X"FD",X"77",X"0C",X"21",X"1B",
		X"8D",X"CD",X"1D",X"94",X"FD",X"73",X"02",X"FD",X"72",X"03",X"C9",X"D6",X"D6",X"EE",X"EE",X"FF",
		X"FF",X"FF",X"FF",X"FD",X"CB",X"01",X"76",X"FD",X"CB",X"01",X"F6",X"FD",X"CB",X"01",X"B6",X"FD",
		X"CB",X"01",X"46",X"28",X"0E",X"1E",X"01",X"3A",X"44",X"48",X"FD",X"BE",X"07",X"30",X"10",X"1E",
		X"04",X"18",X"0C",X"1E",X"02",X"3A",X"42",X"48",X"FD",X"BE",X"05",X"38",X"02",X"1E",X"08",X"D5",
		X"CD",X"C4",X"8E",X"D1",X"A3",X"5F",X"D5",X"CD",X"B5",X"8D",X"D1",X"A3",X"5F",X"D5",X"CD",X"94",
		X"8D",X"D1",X"A3",X"C2",X"44",X"8B",X"CD",X"C4",X"8E",X"5F",X"C3",X"B3",X"8C",X"FD",X"66",X"05",
		X"FD",X"6E",X"07",X"CD",X"1E",X"92",X"01",X"00",X"04",X"E5",X"F5",X"CD",X"D4",X"8D",X"F1",X"E1",
		X"3E",X"02",X"BB",X"28",X"08",X"3E",X"03",X"BB",X"28",X"03",X"B7",X"18",X"01",X"3F",X"CB",X"11",
		X"10",X"E7",X"79",X"C9",X"FD",X"66",X"05",X"FD",X"6E",X"07",X"CD",X"1E",X"92",X"3E",X"04",X"01",
		X"00",X"04",X"E5",X"F5",X"CD",X"D4",X"8D",X"F1",X"E1",X"BB",X"CB",X"11",X"10",X"F4",X"79",X"B7",
		X"C0",X"3E",X"01",X"18",X"EA",X"FD",X"66",X"05",X"FD",X"6E",X"07",X"CD",X"1E",X"92",X"01",X"00",
		X"04",X"C5",X"E5",X"CD",X"D4",X"8D",X"E1",X"7B",X"FE",X"14",X"28",X"01",X"37",X"C1",X"CB",X"11",
		X"10",X"EF",X"79",X"C9",X"E5",X"78",X"21",X"F1",X"8D",X"3D",X"CD",X"1D",X"94",X"E1",X"19",X"7C",
		X"E6",X"03",X"F6",X"44",X"67",X"7D",X"E6",X"1F",X"FE",X"1C",X"38",X"03",X"21",X"00",X"44",X"5E",
		X"C9",X"03",X"00",X"61",X"00",X"1E",X"00",X"C0",X"FF",X"03",X"00",X"30",X"10",X"01",X"10",X"00",
		X"10",X"03",X"00",X"00",X"10",X"01",X"10",X"30",X"10",X"21",X"39",X"8E",X"18",X"03",X"21",X"25",
		X"8E",X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",X"3D",X"CD",X"1D",X"94",X"FD",X"73",
		X"02",X"FD",X"72",X"03",X"C9",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",
		X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"D6",X"6D",X"DB",X"EE",X"EE",X"D6",
		X"D6",X"EE",X"EE",X"EE",X"EE",X"D6",X"D6",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"3A",X"24",X"4A",
		X"FE",X"02",X"38",X"02",X"3E",X"02",X"21",X"6B",X"8E",X"CD",X"1D",X"94",X"EB",X"ED",X"5F",X"E6",
		X"03",X"CD",X"1D",X"94",X"FD",X"73",X"0A",X"FD",X"72",X"0B",X"C9",X"71",X"8E",X"79",X"8E",X"81",
		X"8E",X"80",X"00",X"50",X"00",X"90",X"00",X"A0",X"00",X"50",X"00",X"60",X"00",X"70",X"00",X"50",
		X"00",X"30",X"00",X"50",X"00",X"20",X"00",X"40",X"00",X"00",X"FF",X"01",X"00",X"00",X"01",X"FF",
		X"00",X"06",X"03",X"3A",X"AA",X"49",X"FE",X"04",X"D8",X"06",X"04",X"C9",X"FD",X"7E",X"09",X"B7",
		X"C2",X"DD",X"88",X"FD",X"6E",X"0A",X"FD",X"66",X"0B",X"7E",X"FD",X"77",X"09",X"23",X"FD",X"7E",
		X"01",X"E6",X"F0",X"B6",X"FD",X"77",X"01",X"23",X"FD",X"75",X"0A",X"FD",X"74",X"0B",X"CD",X"44",
		X"8B",X"C3",X"DD",X"88",X"01",X"00",X"04",X"C5",X"21",X"F0",X"8E",X"05",X"78",X"CD",X"17",X"94",
		X"4E",X"23",X"46",X"FD",X"66",X"05",X"FD",X"6E",X"07",X"CD",X"A5",X"91",X"3A",X"42",X"48",X"BC",
		X"20",X"06",X"3A",X"44",X"48",X"BD",X"28",X"01",X"37",X"C1",X"CB",X"11",X"10",X"D9",X"79",X"C9",
		X"00",X"F0",X"10",X"00",X"00",X"10",X"F0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"1E",X"00",X"73",X"23",X"0B",X"79",X"B0",X"20",X"F9",X"C9",X"DD",X"46",X"00",X"DD",X"23",X"DD",
		X"4E",X"00",X"AF",X"B9",X"C8",X"DD",X"6E",X"01",X"DD",X"66",X"02",X"DD",X"7E",X"03",X"D5",X"11",
		X"04",X"00",X"DD",X"19",X"D1",X"B7",X"20",X"1F",X"DD",X"5E",X"00",X"DD",X"23",X"B8",X"20",X"08",
		X"C5",X"41",X"CD",X"7D",X"8F",X"C1",X"18",X"D7",X"3E",X"23",X"FF",X"C5",X"06",X"01",X"CD",X"7D",
		X"8F",X"C1",X"0D",X"20",X"F3",X"18",X"C8",X"AF",X"B8",X"20",X"11",X"41",X"C5",X"DD",X"5E",X"00",
		X"DD",X"23",X"06",X"01",X"CD",X"7D",X"8F",X"C1",X"10",X"F2",X"18",X"B3",X"3E",X"23",X"FF",X"C5",
		X"DD",X"5E",X"00",X"DD",X"23",X"06",X"01",X"CD",X"7D",X"8F",X"C1",X"0D",X"20",X"EE",X"18",X"9F",
		X"DD",X"7E",X"00",X"77",X"CD",X"6F",X"90",X"23",X"DD",X"23",X"10",X"F4",X"C9",X"DD",X"7E",X"00",
		X"77",X"CD",X"6F",X"90",X"CD",X"79",X"90",X"DD",X"23",X"10",X"F2",X"C9",X"DD",X"7E",X"00",X"DD",
		X"23",X"B7",X"C8",X"CB",X"7F",X"20",X"25",X"4F",X"DD",X"46",X"00",X"DD",X"23",X"CB",X"78",X"CB",
		X"B8",X"28",X"08",X"23",X"0D",X"28",X"1B",X"10",X"FA",X"18",X"ED",X"DD",X"7E",X"00",X"DD",X"23",
		X"77",X"CD",X"6F",X"90",X"23",X"0D",X"28",X"0A",X"10",X"F6",X"18",X"DC",X"D5",X"CB",X"BF",X"47",
		X"18",X"03",X"D5",X"06",X"01",X"11",X"20",X"00",X"7D",X"E6",X"E0",X"6F",X"19",X"10",X"FD",X"D1",
		X"18",X"BA",X"06",X"01",X"CD",X"80",X"8F",X"DD",X"2B",X"C9",X"0E",X"00",X"1A",X"81",X"0E",X"00",
		X"86",X"FE",X"0A",X"FA",X"E9",X"8F",X"0C",X"D6",X"0A",X"12",X"2B",X"1B",X"10",X"EE",X"C9",X"0E",
		X"00",X"1A",X"91",X"F2",X"FA",X"8F",X"3E",X"09",X"18",X"02",X"0E",X"00",X"96",X"F2",X"04",X"90",
		X"0E",X"01",X"C6",X"0A",X"12",X"2B",X"1B",X"10",X"E8",X"C9",X"AF",X"5F",X"E5",X"C5",X"77",X"CD",
		X"6F",X"90",X"23",X"10",X"F9",X"C1",X"E1",X"CD",X"79",X"90",X"0D",X"20",X"EF",X"C9",X"DD",X"7E",
		X"00",X"05",X"28",X"08",X"FE",X"00",X"20",X"03",X"B9",X"28",X"03",X"0D",X"F6",X"30",X"C5",X"D5",
		X"CD",X"D2",X"8F",X"D1",X"C1",X"DD",X"23",X"78",X"B7",X"20",X"E3",X"C9",X"C5",X"E5",X"CD",X"70",
		X"8F",X"E1",X"CD",X"79",X"90",X"C1",X"0D",X"20",X"F3",X"C9",X"C5",X"E5",X"77",X"CD",X"6F",X"90",
		X"23",X"10",X"F9",X"E1",X"CD",X"79",X"90",X"C1",X"0D",X"20",X"EF",X"C9",X"C5",X"E5",X"77",X"CD",
		X"6F",X"90",X"3C",X"23",X"10",X"F8",X"E1",X"CD",X"79",X"90",X"C1",X"0D",X"20",X"EE",X"C9",X"F5",
		X"E5",X"7C",X"C6",X"04",X"67",X"73",X"E1",X"F1",X"C9",X"D5",X"11",X"20",X"00",X"19",X"D1",X"C9",
		X"1A",X"BE",X"38",X"0B",X"20",X"06",X"13",X"23",X"10",X"F6",X"AF",X"C9",X"3E",X"02",X"C9",X"3E",
		X"01",X"C9",X"E5",X"06",X"06",X"11",X"8D",X"49",X"CD",X"DA",X"8F",X"21",X"BD",X"41",X"06",X"06",
		X"0E",X"00",X"1E",X"04",X"DD",X"21",X"88",X"49",X"CD",X"1E",X"90",X"E1",X"11",X"19",X"48",X"01",
		X"14",X"48",X"3A",X"01",X"48",X"CB",X"6F",X"20",X"06",X"11",X"13",X"48",X"01",X"0E",X"48",X"CB",
		X"7F",X"C8",X"C5",X"F5",X"06",X"06",X"CD",X"DA",X"8F",X"F1",X"DD",X"21",X"0E",X"48",X"21",X"BF",
		X"40",X"CB",X"6F",X"28",X"07",X"DD",X"21",X"14",X"48",X"21",X"FF",X"42",X"06",X"06",X"1E",X"05",
		X"CD",X"1E",X"90",X"E1",X"3A",X"A6",X"49",X"E6",X"0F",X"FE",X"04",X"D0",X"3A",X"80",X"50",X"2F",
		X"E6",X"0C",X"C8",X"CB",X"3F",X"CB",X"3F",X"E5",X"21",X"22",X"91",X"3D",X"CD",X"1D",X"94",X"EB",
		X"3A",X"A6",X"49",X"E6",X"0F",X"CD",X"10",X"94",X"EB",X"E1",X"06",X"06",X"CD",X"80",X"90",X"FE",
		X"02",X"20",X"01",X"C9",X"21",X"A6",X"49",X"34",X"21",X"A7",X"49",X"7E",X"34",X"47",X"CD",X"70",
		X"91",X"C9",X"28",X"91",X"40",X"91",X"58",X"91",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"02",X"05",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"01",X"05",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",
		X"21",X"7C",X"40",X"1E",X"01",X"0E",X"06",X"AF",X"B0",X"28",X"0D",X"3E",X"2D",X"C5",X"CD",X"D2",
		X"8F",X"C1",X"0D",X"10",X"F8",X"AF",X"B9",X"C8",X"41",X"C5",X"CD",X"D2",X"8F",X"C1",X"10",X"F9",
		X"C9",X"7E",X"FE",X"FF",X"C8",X"FF",X"23",X"18",X"F8",X"7E",X"FE",X"FF",X"C8",X"23",X"4E",X"23",
		X"46",X"23",X"FF",X"18",X"F4",X"7D",X"80",X"6F",X"7C",X"81",X"67",X"C9",X"7C",X"FE",X"30",X"38",
		X"36",X"FE",X"E1",X"30",X"32",X"06",X"0C",X"1E",X"84",X"3E",X"D0",X"BC",X"38",X"0A",X"D6",X"10",
		X"57",X"7B",X"D6",X"0C",X"5F",X"7A",X"10",X"F3",X"7D",X"FE",X"40",X"38",X"1A",X"FE",X"F1",X"30",
		X"16",X"06",X"0C",X"3E",X"EF",X"BD",X"38",X"07",X"1C",X"D6",X"10",X"10",X"F8",X"1E",X"00",X"21",
		X"68",X"48",X"16",X"00",X"19",X"7E",X"C9",X"3E",X"FF",X"C9",X"B7",X"06",X"08",X"26",X"00",X"6F",
		X"1E",X"0C",X"ED",X"6A",X"7C",X"38",X"03",X"BB",X"38",X"03",X"93",X"67",X"AF",X"3F",X"10",X"F2",
		X"CB",X"15",X"CB",X"25",X"CB",X"25",X"CB",X"25",X"CB",X"25",X"7D",X"C6",X"30",X"6C",X"67",X"CB",
		X"25",X"CB",X"25",X"CB",X"25",X"CB",X"25",X"3E",X"10",X"85",X"ED",X"44",X"6F",X"C9",X"7D",X"ED",
		X"44",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"5F",X"3E",X"F0",X"84",X"E6",X"F8",X"26",X"00",X"6F",
		X"29",X"29",X"16",X"40",X"19",X"C9",X"21",X"68",X"48",X"01",X"90",X"00",X"CD",X"00",X"8F",X"3A",
		X"AA",X"49",X"FE",X"05",X"30",X"18",X"3D",X"21",X"F5",X"93",X"CD",X"1D",X"94",X"21",X"68",X"48",
		X"1A",X"13",X"FE",X"FF",X"28",X"08",X"06",X"00",X"4F",X"09",X"36",X"20",X"18",X"EF",X"21",X"30",
		X"93",X"3A",X"AA",X"49",X"FE",X"07",X"38",X"02",X"3E",X"07",X"3D",X"16",X"00",X"5F",X"19",X"46",
		X"C5",X"CD",X"F0",X"92",X"C1",X"10",X"F9",X"3A",X"AA",X"49",X"FE",X"0A",X"38",X"02",X"3E",X"0A",
		X"3D",X"21",X"37",X"93",X"CD",X"1D",X"94",X"EB",X"7E",X"B7",X"C2",X"AA",X"92",X"21",X"AA",X"48",
		X"7E",X"E6",X"F0",X"28",X"0E",X"E5",X"23",X"7E",X"E6",X"F0",X"20",X"FA",X"D1",X"EB",X"4E",X"1A",
		X"77",X"79",X"12",X"7E",X"E6",X"0F",X"F6",X"30",X"77",X"C9",X"4F",X"23",X"46",X"23",X"E5",X"21",
		X"68",X"48",X"ED",X"5F",X"E6",X"7F",X"CB",X"27",X"5F",X"ED",X"5F",X"E6",X"3F",X"83",X"5F",X"16",
		X"00",X"19",X"B7",X"E5",X"11",X"F8",X"48",X"ED",X"52",X"EB",X"E1",X"38",X"04",X"21",X"68",X"48",
		X"19",X"7E",X"B7",X"28",X"15",X"23",X"23",X"23",X"23",X"23",X"E5",X"11",X"F8",X"48",X"ED",X"52",
		X"E1",X"38",X"EE",X"11",X"90",X"00",X"ED",X"52",X"18",X"E7",X"71",X"10",X"C2",X"E1",X"18",X"98",
		X"21",X"82",X"48",X"ED",X"5F",X"5F",X"ED",X"5F",X"83",X"5F",X"ED",X"5F",X"E6",X"07",X"B7",X"28",
		X"05",X"3D",X"CB",X"03",X"18",X"F8",X"7B",X"E6",X"07",X"5F",X"ED",X"5F",X"57",X"ED",X"5F",X"E6",
		X"0F",X"B7",X"28",X"05",X"3D",X"CB",X"02",X"18",X"F8",X"7A",X"E6",X"07",X"16",X"00",X"19",X"B7",
		X"28",X"07",X"3D",X"11",X"0C",X"00",X"19",X"18",X"F6",X"AF",X"BE",X"20",X"C3",X"36",X"40",X"C9",
		X"01",X"02",X"03",X"04",X"05",X"06",X"07",X"4B",X"93",X"5C",X"93",X"6D",X"93",X"7E",X"93",X"8F",
		X"93",X"A0",X"93",X"B1",X"93",X"C2",X"93",X"D3",X"93",X"E4",X"93",X"11",X"03",X"12",X"03",X"13",
		X"03",X"14",X"03",X"01",X"0F",X"02",X"1E",X"04",X"2E",X"03",X"24",X"00",X"11",X"03",X"12",X"03",
		X"13",X"03",X"14",X"04",X"01",X"0F",X"02",X"1D",X"04",X"31",X"03",X"21",X"00",X"11",X"02",X"12",
		X"02",X"13",X"04",X"14",X"04",X"01",X"0E",X"02",X"20",X"04",X"2F",X"03",X"22",X"00",X"11",X"02",
		X"12",X"02",X"13",X"04",X"14",X"05",X"01",X"0E",X"02",X"1E",X"04",X"2F",X"03",X"23",X"00",X"11",
		X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1C",X"04",X"31",X"03",X"24",X"00",
		X"11",X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1B",X"04",X"31",X"03",X"24",
		X"00",X"11",X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1C",X"04",X"31",X"03",
		X"22",X"00",X"11",X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1C",X"04",X"31",
		X"03",X"22",X"00",X"11",X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1C",X"04",
		X"31",X"03",X"22",X"00",X"11",X"02",X"12",X"02",X"13",X"05",X"14",X"05",X"01",X"0C",X"02",X"1C",
		X"04",X"31",X"03",X"22",X"00",X"FD",X"93",X"02",X"94",X"06",X"94",X"09",X"94",X"1E",X"3E",X"45",
		X"72",X"FF",X"1E",X"3E",X"72",X"FF",X"3E",X"72",X"FF",X"3E",X"FF",X"5F",X"87",X"83",X"18",X"08",
		X"87",X"5F",X"87",X"83",X"18",X"02",X"87",X"87",X"16",X"00",X"5F",X"19",X"C9",X"CD",X"17",X"94",
		X"5E",X"23",X"56",X"C9",X"06",X"04",X"0E",X"00",X"CB",X"3F",X"38",X"03",X"0C",X"10",X"F9",X"79",
		X"C9",X"0E",X"01",X"B7",X"28",X"05",X"3D",X"CB",X"21",X"18",X"F8",X"79",X"C9",X"DD",X"21",X"82",
		X"40",X"01",X"0C",X"0C",X"FD",X"21",X"68",X"48",X"C5",X"DD",X"E5",X"C5",X"21",X"75",X"94",X"FD",
		X"7E",X"00",X"CB",X"9F",X"FD",X"77",X"00",X"CB",X"7F",X"20",X"03",X"21",X"7F",X"94",X"4F",X"E6",
		X"70",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CD",X"1D",X"94",X"EB",X"11",X"93",X"94",
		X"D5",X"79",X"E6",X"07",X"E9",X"AD",X"94",X"AD",X"94",X"B2",X"94",X"AD",X"94",X"B2",X"94",X"C0",
		X"94",X"C0",X"94",X"B2",X"94",X"C0",X"94",X"C0",X"94",X"A8",X"94",X"A8",X"94",X"B2",X"94",X"B6",
		X"2D",X"B9",X"94",X"FD",X"23",X"DD",X"23",X"DD",X"23",X"C1",X"10",X"AF",X"DD",X"E1",X"01",X"40",
		X"00",X"DD",X"09",X"C1",X"0D",X"20",X"A1",X"C9",X"CD",X"76",X"95",X"18",X"20",X"CD",X"87",X"95",
		X"18",X"1B",X"3E",X"88",X"1E",X"14",X"C3",X"CD",X"94",X"3E",X"01",X"1E",X"0A",X"C3",X"CD",X"94",
		X"AF",X"1E",X"16",X"01",X"02",X"02",X"DD",X"E5",X"E1",X"CD",X"4A",X"90",X"C9",X"DD",X"E5",X"E1",
		X"01",X"02",X"02",X"CD",X"5C",X"90",X"C9",X"06",X"04",X"C5",X"CD",X"2D",X"95",X"3E",X"23",X"06",
		X"1E",X"FF",X"06",X"90",X"21",X"68",X"48",X"C5",X"E5",X"7E",X"F5",X"B7",X"11",X"68",X"48",X"ED",
		X"52",X"7D",X"CD",X"EA",X"91",X"CD",X"1E",X"92",X"F1",X"FE",X"20",X"20",X"0C",X"3E",X"88",X"1E",
		X"14",X"01",X"02",X"02",X"CD",X"5C",X"90",X"18",X"14",X"E6",X"70",X"FE",X"30",X"20",X"05",X"CD",
		X"B6",X"2D",X"18",X"09",X"AF",X"1E",X"16",X"01",X"02",X"02",X"CD",X"0C",X"90",X"E1",X"23",X"C1",
		X"10",X"C5",X"3E",X"23",X"06",X"3C",X"FF",X"C1",X"05",X"C2",X"D9",X"94",X"C9",X"FD",X"21",X"68",
		X"48",X"01",X"0C",X"0C",X"DD",X"21",X"82",X"40",X"C5",X"DD",X"E5",X"C5",X"21",X"75",X"94",X"FD",
		X"7E",X"00",X"CB",X"7F",X"20",X"03",X"21",X"89",X"94",X"4F",X"E6",X"70",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CD",X"1D",X"94",X"EB",X"11",X"60",X"95",X"D5",X"79",X"E6",X"07",X"E9",
		X"FD",X"23",X"DD",X"23",X"DD",X"23",X"C1",X"10",X"D2",X"DD",X"E1",X"11",X"40",X"00",X"DD",X"19",
		X"C1",X"0D",X"C2",X"38",X"95",X"C9",X"21",X"7F",X"95",X"3D",X"CD",X"1D",X"94",X"7A",X"C9",X"0D",
		X"C0",X"0E",X"C4",X"0F",X"C8",X"10",X"CC",X"F5",X"3A",X"01",X"48",X"CB",X"7F",X"20",X"04",X"3E",
		X"07",X"18",X"03",X"3A",X"AA",X"49",X"FE",X"08",X"38",X"04",X"D6",X"07",X"18",X"F8",X"21",X"B3",
		X"95",X"3D",X"16",X"00",X"5F",X"19",X"4E",X"21",X"BA",X"95",X"F1",X"3D",X"16",X"00",X"5F",X"19",
		X"5E",X"79",X"C9",X"D8",X"E0",X"E4",X"D4",X"E8",X"EC",X"DC",X"06",X"07",X"08",X"09",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"20",X"4F",X"21",X"45",X"48",X"06",X"1E",X"CF",X"21",X"20",X"4A",X"06",X"56",X"CF",X"CD",
		X"3A",X"97",X"C5",X"3A",X"AB",X"49",X"32",X"20",X"4A",X"FE",X"04",X"30",X"0D",X"ED",X"5F",X"E6",
		X"03",X"FE",X"03",X"38",X"02",X"3E",X"02",X"32",X"21",X"4A",X"21",X"70",X"97",X"CD",X"4D",X"97",
		X"FD",X"21",X"26",X"4A",X"C5",X"FD",X"E5",X"D1",X"01",X"04",X"00",X"ED",X"B0",X"11",X"0E",X"00",
		X"FD",X"19",X"C1",X"10",X"EF",X"C1",X"C5",X"21",X"7E",X"98",X"CD",X"4D",X"97",X"FD",X"21",X"22",
		X"4A",X"5E",X"23",X"56",X"23",X"FD",X"73",X"02",X"FD",X"72",X"03",X"11",X"0E",X"00",X"FD",X"19",
		X"10",X"EF",X"C1",X"21",X"2C",X"99",X"CD",X"4D",X"97",X"FD",X"21",X"22",X"4A",X"5E",X"23",X"56",
		X"23",X"FD",X"73",X"0A",X"FD",X"73",X"0C",X"FD",X"72",X"0B",X"FD",X"72",X"0D",X"11",X"0E",X"00",
		X"FD",X"19",X"10",X"E9",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",X"22",X"4A",X"DD",X"21",X"45",
		X"48",X"CD",X"3A",X"97",X"C5",X"FD",X"36",X"00",X"03",X"FD",X"7E",X"08",X"B7",X"20",X"07",X"FD",
		X"36",X"08",X"05",X"CD",X"29",X"89",X"FD",X"35",X"08",X"FD",X"7E",X"09",X"B7",X"C2",X"FC",X"96",
		X"FD",X"6E",X"0C",X"FD",X"66",X"0D",X"7E",X"FE",X"FF",X"20",X"0F",X"3A",X"AB",X"49",X"FE",X"06",
		X"CA",X"E7",X"96",X"FD",X"6E",X"0A",X"FD",X"66",X"0B",X"7E",X"23",X"5E",X"23",X"FD",X"75",X"0C",
		X"FD",X"74",X"0D",X"FD",X"77",X"01",X"FD",X"73",X"09",X"21",X"F8",X"96",X"16",X"00",X"5F",X"19",
		X"7E",X"FD",X"77",X"04",X"C3",X"FC",X"96",X"FD",X"7E",X"07",X"21",X"23",X"9C",X"FE",X"80",X"D2",
		X"C9",X"96",X"21",X"CC",X"9B",X"C3",X"C9",X"96",X"2B",X"A8",X"2B",X"28",X"CD",X"19",X"8B",X"D2",
		X"08",X"97",X"CD",X"DD",X"88",X"C3",X"08",X"97",X"DD",X"E5",X"D1",X"13",X"FD",X"E5",X"E1",X"23",
		X"23",X"23",X"23",X"01",X"04",X"00",X"ED",X"B0",X"DD",X"36",X"00",X"00",X"11",X"0E",X"00",X"FD",
		X"19",X"11",X"05",X"00",X"DD",X"19",X"C1",X"05",X"C2",X"94",X"96",X"3A",X"20",X"4A",X"B7",X"20",
		X"02",X"ED",X"5F",X"3D",X"32",X"20",X"4A",X"C3",X"84",X"96",X"3A",X"AB",X"49",X"21",X"46",X"97",
		X"16",X"00",X"5F",X"19",X"46",X"C9",X"05",X"05",X"05",X"05",X"06",X"06",X"06",X"3A",X"20",X"4A",
		X"CD",X"1D",X"94",X"EB",X"FE",X"08",X"D0",X"3A",X"21",X"4A",X"CD",X"1D",X"94",X"EB",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7E",X"97",X"84",X"97",X"8A",X"97",X"90",X"97",X"36",X"98",X"4E",X"98",X"66",X"98",X"96",X"97",
		X"AA",X"97",X"AA",X"97",X"BE",X"97",X"D2",X"97",X"D2",X"97",X"E6",X"97",X"FA",X"97",X"FA",X"97",
		X"0E",X"98",X"22",X"98",X"22",X"98",X"28",X"B0",X"52",X"E0",X"2B",X"40",X"52",X"D0",X"A8",X"90",
		X"52",X"98",X"A8",X"60",X"52",X"B0",X"28",X"A0",X"52",X"60",X"2B",X"B0",X"52",X"E0",X"28",X"40",
		X"52",X"D0",X"28",X"90",X"52",X"98",X"2B",X"60",X"52",X"B0",X"2B",X"A0",X"52",X"60",X"2B",X"B0",
		X"52",X"98",X"28",X"80",X"52",X"E0",X"A8",X"50",X"52",X"98",X"A8",X"80",X"52",X"60",X"2B",X"A0",
		X"52",X"B8",X"28",X"B0",X"52",X"98",X"A8",X"80",X"52",X"E0",X"2B",X"50",X"52",X"98",X"A8",X"80",
		X"52",X"60",X"28",X"A0",X"52",X"B8",X"2B",X"C0",X"52",X"98",X"28",X"A0",X"52",X"E0",X"2B",X"90",
		X"52",X"D0",X"2B",X"60",X"52",X"B0",X"A8",X"80",X"52",X"60",X"28",X"C0",X"52",X"98",X"A8",X"A0",
		X"52",X"E0",X"28",X"90",X"52",X"D0",X"A8",X"60",X"52",X"B0",X"28",X"80",X"52",X"60",X"28",X"A0",
		X"52",X"E0",X"2B",X"A0",X"52",X"A0",X"A8",X"40",X"52",X"C0",X"28",X"80",X"52",X"70",X"2B",X"A0",
		X"52",X"60",X"2B",X"A0",X"52",X"E0",X"28",X"A0",X"52",X"A0",X"2B",X"40",X"52",X"C0",X"2B",X"80",
		X"52",X"70",X"28",X"A0",X"52",X"60",X"A8",X"50",X"52",X"E0",X"28",X"E0",X"52",X"C8",X"28",X"80",
		X"52",X"B0",X"28",X"A0",X"52",X"90",X"A8",X"50",X"52",X"78",X"A8",X"40",X"52",X"60",X"28",X"E0",
		X"52",X"D8",X"A8",X"60",X"52",X"C0",X"28",X"B0",X"52",X"A8",X"A8",X"40",X"52",X"90",X"28",X"90",
		X"52",X"78",X"A8",X"50",X"52",X"60",X"28",X"A0",X"52",X"48",X"A8",X"30",X"52",X"70",X"28",X"88",
		X"52",X"88",X"A8",X"50",X"52",X"A8",X"28",X"E8",X"52",X"C0",X"28",X"D0",X"52",X"F0",X"8C",X"98",
		X"92",X"98",X"98",X"98",X"9E",X"98",X"08",X"99",X"14",X"99",X"20",X"99",X"A4",X"98",X"AE",X"98",
		X"B8",X"98",X"C2",X"98",X"CC",X"98",X"D6",X"98",X"E0",X"98",X"E0",X"98",X"EA",X"98",X"F4",X"98",
		X"F4",X"98",X"FE",X"98",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"D6",X"D6",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",X"FF",X"FF",
		X"FF",X"FF",X"EE",X"EE",X"FF",X"FF",X"D6",X"D6",X"EE",X"EE",X"AA",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"D6",X"D6",X"FF",X"FF",X"AA",X"AA",X"EE",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"D6",X"D6",X"FF",X"FF",X"D6",X"D6",X"AA",X"AA",X"FF",X"FF",X"AA",X"AA",X"EE",X"EE",
		X"AA",X"AA",X"AA",X"AA",X"AA",X"AA",X"EE",X"EE",X"AA",X"AA",X"D6",X"D6",X"3A",X"99",X"40",X"99",
		X"46",X"99",X"4C",X"99",X"4E",X"9B",X"7E",X"9B",X"C0",X"9B",X"52",X"99",X"5C",X"99",X"5C",X"99",
		X"F4",X"99",X"FE",X"99",X"FE",X"99",X"6A",X"9A",X"74",X"9A",X"74",X"9A",X"E0",X"9A",X"EA",X"9A",
		X"EA",X"9A",X"66",X"99",X"77",X"99",X"88",X"99",X"9B",X"99",X"A4",X"99",X"AD",X"99",X"BE",X"99",
		X"CF",X"99",X"E2",X"99",X"EB",X"99",X"03",X"60",X"00",X"10",X"03",X"10",X"00",X"38",X"01",X"80",
		X"02",X"38",X"03",X"10",X"02",X"10",X"FF",X"00",X"38",X"01",X"80",X"02",X"38",X"03",X"10",X"02",
		X"10",X"03",X"60",X"00",X"10",X"03",X"10",X"FF",X"01",X"30",X"02",X"38",X"03",X"10",X"02",X"10",
		X"03",X"60",X"00",X"10",X"03",X"10",X"00",X"38",X"01",X"50",X"FF",X"01",X"40",X"00",X"50",X"03",
		X"40",X"02",X"50",X"FF",X"03",X"40",X"02",X"50",X"01",X"40",X"00",X"50",X"FF",X"00",X"10",X"01",
		X"10",X"00",X"38",X"03",X"80",X"02",X"38",X"01",X"10",X"02",X"10",X"01",X"60",X"FF",X"01",X"10",
		X"02",X"10",X"01",X"60",X"00",X"10",X"01",X"10",X"00",X"38",X"03",X"80",X"02",X"38",X"FF",X"03",
		X"50",X"02",X"38",X"01",X"10",X"02",X"10",X"01",X"60",X"00",X"10",X"01",X"10",X"00",X"38",X"03",
		X"30",X"FF",X"00",X"50",X"01",X"40",X"02",X"50",X"03",X"40",X"FF",X"02",X"50",X"03",X"40",X"00",
		X"50",X"01",X"40",X"FF",X"08",X"9A",X"11",X"9A",X"1C",X"9A",X"25",X"9A",X"30",X"9A",X"39",X"9A",
		X"42",X"9A",X"4D",X"9A",X"56",X"9A",X"61",X"9A",X"02",X"48",X"03",X"60",X"00",X"48",X"01",X"60",
		X"FF",X"03",X"30",X"00",X"48",X"01",X"60",X"02",X"48",X"03",X"30",X"FF",X"01",X"60",X"02",X"48",
		X"03",X"60",X"00",X"48",X"FF",X"03",X"20",X"02",X"58",X"01",X"40",X"00",X"58",X"03",X"20",X"FF",
		X"00",X"58",X"03",X"40",X"02",X"58",X"01",X"40",X"FF",X"03",X"60",X"02",X"48",X"01",X"60",X"00",
		X"48",X"FF",X"01",X"30",X"00",X"48",X"03",X"60",X"02",X"48",X"01",X"30",X"FF",X"02",X"48",X"01",
		X"60",X"00",X"48",X"03",X"60",X"FF",X"01",X"20",X"02",X"58",X"03",X"40",X"00",X"58",X"01",X"20",
		X"FF",X"03",X"40",X"00",X"58",X"01",X"40",X"02",X"58",X"FF",X"7E",X"9A",X"87",X"9A",X"92",X"9A",
		X"9B",X"9A",X"A4",X"9A",X"AF",X"9A",X"B8",X"9A",X"C3",X"9A",X"CC",X"9A",X"D5",X"9A",X"02",X"48",
		X"03",X"50",X"00",X"48",X"01",X"50",X"FF",X"03",X"30",X"00",X"48",X"01",X"50",X"02",X"48",X"03",
		X"20",X"FF",X"00",X"38",X"03",X"50",X"02",X"38",X"01",X"50",X"FF",X"00",X"40",X"01",X"40",X"02",
		X"40",X"03",X"40",X"FF",X"01",X"10",X"02",X"20",X"03",X"20",X"00",X"20",X"01",X"10",X"FF",X"03",
		X"50",X"02",X"48",X"01",X"50",X"00",X"48",X"FF",X"01",X"20",X"00",X"48",X"03",X"50",X"02",X"48",
		X"01",X"30",X"FF",X"03",X"50",X"00",X"38",X"01",X"50",X"02",X"38",X"FF",X"01",X"40",X"00",X"40",
		X"03",X"40",X"02",X"40",X"FF",X"03",X"10",X"02",X"20",X"01",X"20",X"00",X"20",X"03",X"10",X"FF",
		X"F4",X"9A",X"FD",X"9A",X"06",X"9B",X"0F",X"9B",X"18",X"9B",X"21",X"9B",X"2A",X"9B",X"33",X"9B",
		X"3C",X"9B",X"45",X"9B",X"03",X"40",X"00",X"20",X"01",X"40",X"02",X"20",X"FF",X"02",X"20",X"03",
		X"20",X"00",X"20",X"01",X"20",X"FF",X"01",X"20",X"00",X"20",X"03",X"20",X"02",X"20",X"FF",X"03",
		X"20",X"02",X"20",X"01",X"20",X"00",X"20",X"FF",X"02",X"20",X"03",X"20",X"00",X"20",X"01",X"20",
		X"FF",X"00",X"20",X"03",X"40",X"02",X"20",X"01",X"40",X"FF",X"03",X"20",X"02",X"20",X"01",X"20",
		X"00",X"20",X"FF",X"00",X"20",X"01",X"20",X"02",X"20",X"03",X"20",X"FF",X"02",X"20",X"03",X"20",
		X"00",X"20",X"01",X"20",X"FF",X"03",X"20",X"02",X"20",X"01",X"20",X"00",X"20",X"FF",X"5A",X"9B",
		X"5F",X"9B",X"64",X"9B",X"6B",X"9B",X"70",X"9B",X"77",X"9B",X"01",X"90",X"03",X"90",X"FF",X"03",
		X"B0",X"01",X"B0",X"FF",X"03",X"50",X"01",X"A0",X"03",X"50",X"FF",X"03",X"70",X"01",X"70",X"FF",
		X"01",X"50",X"03",X"70",X"01",X"20",X"FF",X"01",X"60",X"03",X"70",X"01",X"10",X"FF",X"8A",X"9B",
		X"93",X"9B",X"9C",X"9B",X"A5",X"9B",X"AE",X"9B",X"B7",X"9B",X"03",X"90",X"02",X"08",X"01",X"90",
		X"00",X"08",X"FF",X"01",X"70",X"02",X"08",X"03",X"70",X"00",X"08",X"FF",X"03",X"60",X"02",X"08",
		X"01",X"60",X"00",X"08",X"FF",X"01",X"60",X"02",X"08",X"03",X"60",X"00",X"08",X"FF",X"03",X"60",
		X"02",X"08",X"01",X"60",X"00",X"08",X"FF",X"01",X"50",X"02",X"08",X"03",X"50",X"00",X"08",X"FF",
		X"CC",X"9B",X"E0",X"9B",X"EC",X"9B",X"47",X"9C",X"3B",X"9C",X"23",X"9C",X"03",X"38",X"02",X"08",
		X"01",X"28",X"02",X"08",X"03",X"50",X"02",X"08",X"01",X"40",X"02",X"08",X"03",X"50",X"02",X"08",
		X"01",X"50",X"02",X"08",X"03",X"60",X"02",X"08",X"01",X"68",X"02",X"08",X"03",X"60",X"02",X"08",
		X"01",X"90",X"02",X"08",X"03",X"78",X"02",X"08",X"01",X"98",X"02",X"08",X"03",X"88",X"02",X"08",
		X"01",X"98",X"02",X"08",X"03",X"90",X"02",X"08",X"01",X"90",X"02",X"08",X"03",X"60",X"02",X"08",
		X"01",X"60",X"02",X"08",X"03",X"68",X"02",X"08",X"01",X"58",X"02",X"08",X"03",X"28",X"02",X"08",
		X"01",X"20",X"FF",X"03",X"20",X"00",X"08",X"01",X"28",X"00",X"08",X"03",X"58",X"00",X"08",X"01",
		X"68",X"00",X"08",X"03",X"60",X"00",X"08",X"01",X"60",X"00",X"08",X"03",X"90",X"00",X"08",X"01",
		X"90",X"00",X"08",X"03",X"98",X"00",X"08",X"01",X"88",X"00",X"08",X"03",X"98",X"00",X"08",X"01",
		X"78",X"00",X"08",X"03",X"90",X"00",X"08",X"01",X"60",X"00",X"08",X"03",X"68",X"00",X"08",X"01",
		X"60",X"00",X"08",X"03",X"50",X"00",X"08",X"01",X"50",X"00",X"08",X"03",X"40",X"00",X"08",X"01",
		X"50",X"00",X"08",X"03",X"28",X"00",X"08",X"01",X"38",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CE",X"9C",X"DA",X"9C",X"1C",X"9D",X"A0",X"9D",X"AD",X"9D",X"AD",X"9D",X"D0",X"9D",X"FB",X"9D",
		X"0A",X"9E",X"18",X"9E",X"63",X"9E",X"63",X"9E",X"7A",X"9E",X"C6",X"9E",X"F6",X"9E",X"05",X"9F",
		X"11",X"9F",X"24",X"9F",X"00",X"A0",X"68",X"A0",X"7E",X"A0",X"96",X"A0",X"1C",X"A1",X"D4",X"A3",
		X"E2",X"A3",X"F9",X"A3",X"07",X"A4",X"25",X"A4",X"5C",X"A4",X"69",X"A4",X"B3",X"A4",X"81",X"01",
		X"01",X"D3",X"9C",X"E8",X"09",X"05",X"40",X"37",X"39",X"FF",X"01",X"00",X"04",X"E4",X"9C",X"82",
		X"00",X"04",X"00",X"9D",X"EA",X"10",X"05",X"51",X"50",X"4B",X"4A",X"49",X"48",X"47",X"46",X"45",
		X"B5",X"40",X"41",X"42",X"43",X"44",X"45",X"46",X"90",X"D4",X"E8",X"21",X"10",X"25",X"B6",X"FF",
		X"EA",X"10",X"05",X"45",X"43",X"41",X"3B",X"39",X"37",X"35",X"33",X"31",X"B5",X"4A",X"50",X"52",
		X"54",X"56",X"58",X"5A",X"90",X"D4",X"E8",X"21",X"10",X"30",X"B6",X"FF",X"01",X"00",X"02",X"26",
		X"9D",X"82",X"00",X"03",X"63",X"9D",X"AD",X"58",X"57",X"56",X"55",X"54",X"53",X"55",X"54",X"53",
		X"52",X"51",X"50",X"52",X"51",X"50",X"49",X"48",X"47",X"49",X"48",X"47",X"46",X"45",X"44",X"46",
		X"45",X"44",X"43",X"42",X"41",X"43",X"42",X"41",X"40",X"39",X"38",X"40",X"39",X"38",X"37",X"36",
		X"35",X"37",X"36",X"35",X"34",X"33",X"32",X"34",X"33",X"32",X"31",X"30",X"29",X"31",X"30",X"29",
		X"28",X"27",X"FF",X"AD",X"55",X"54",X"53",X"52",X"51",X"50",X"52",X"51",X"50",X"4B",X"4A",X"50",
		X"4B",X"4A",X"49",X"48",X"47",X"46",X"48",X"47",X"46",X"45",X"44",X"46",X"45",X"44",X"43",X"42",
		X"44",X"43",X"42",X"41",X"40",X"42",X"41",X"40",X"3B",X"3A",X"39",X"3B",X"3A",X"39",X"38",X"37",
		X"39",X"E9",X"07",X"30",X"C0",X"07",X"59",X"5A",X"5B",X"60",X"61",X"62",X"63",X"64",X"65",X"FF",
		X"C1",X"01",X"03",X"A5",X"9D",X"E8",X"06",X"06",X"C0",X"40",X"0F",X"D1",X"FF",X"82",X"00",X"03",
		X"B2",X"9D",X"E8",X"18",X"10",X"C0",X"1F",X"10",X"B6",X"C1",X"AF",X"19",X"14",X"18",X"12",X"17",
		X"1A",X"14",X"17",X"1A",X"15",X"21",X"19",X"15",X"18",X"1B",X"16",X"19",X"14",X"17",X"1B",X"FF",
		X"82",X"00",X"05",X"D5",X"9D",X"AD",X"C0",X"1F",X"39",X"4A",X"4B",X"50",X"51",X"52",X"53",X"54",
		X"B5",X"50",X"4B",X"4A",X"39",X"38",X"37",X"36",X"35",X"34",X"33",X"32",X"31",X"30",X"2B",X"2A",
		X"29",X"28",X"27",X"26",X"25",X"24",X"23",X"22",X"21",X"20",X"FF",X"84",X"01",X"03",X"00",X"9E",
		X"E8",X"04",X"06",X"34",X"50",X"45",X"42",X"36",X"32",X"FF",X"84",X"00",X"03",X"0F",X"9E",X"B3",
		X"E8",X"05",X"01",X"C0",X"28",X"50",X"B9",X"FF",X"01",X"00",X"04",X"27",X"9E",X"02",X"00",X"04",
		X"3B",X"9E",X"84",X"00",X"04",X"4F",X"9E",X"AD",X"40",X"B3",X"50",X"B3",X"4B",X"B3",X"49",X"B3",
		X"47",X"B3",X"45",X"B3",X"44",X"B3",X"42",X"B3",X"40",X"B6",X"FF",X"AD",X"37",X"B3",X"47",X"B3",
		X"45",X"B3",X"44",X"B3",X"42",X"B3",X"40",X"B3",X"3B",X"B3",X"39",X"B3",X"37",X"B6",X"FF",X"AD",
		X"34",X"B3",X"44",X"B3",X"42",X"B3",X"40",X"B3",X"3B",X"B3",X"39",X"B3",X"37",X"B3",X"35",X"B3",
		X"34",X"B6",X"FF",X"82",X"00",X"03",X"68",X"9E",X"E8",X"05",X"09",X"3B",X"3A",X"39",X"38",X"37",
		X"36",X"B5",X"35",X"34",X"33",X"32",X"31",X"30",X"B3",X"FF",X"82",X"00",X"02",X"7F",X"9E",X"AD",
		X"58",X"57",X"56",X"55",X"54",X"53",X"55",X"54",X"53",X"52",X"51",X"50",X"52",X"51",X"50",X"49",
		X"48",X"47",X"49",X"48",X"47",X"46",X"45",X"44",X"46",X"45",X"44",X"43",X"42",X"41",X"43",X"42",
		X"41",X"40",X"39",X"38",X"40",X"39",X"38",X"37",X"36",X"35",X"37",X"36",X"35",X"34",X"33",X"32",
		X"34",X"33",X"32",X"31",X"30",X"29",X"31",X"30",X"29",X"28",X"27",X"FF",X"40",X"B7",X"D1",X"40",
		X"B7",X"D1",X"40",X"B7",X"D9",X"FF",X"01",X"00",X"05",X"D5",X"9E",X"02",X"00",X"05",X"E0",X"9E",
		X"84",X"00",X"05",X"EB",X"9E",X"E9",X"10",X"20",X"5B",X"50",X"53",X"58",X"BF",X"56",X"57",X"FF",
		X"E9",X"10",X"20",X"46",X"42",X"48",X"45",X"BF",X"40",X"49",X"FF",X"E9",X"10",X"20",X"60",X"68",
		X"63",X"66",X"BF",X"69",X"67",X"FF",X"81",X"01",X"03",X"FB",X"9E",X"E8",X"10",X"10",X"54",X"50",
		X"54",X"50",X"54",X"50",X"FF",X"81",X"01",X"01",X"0A",X"9F",X"E8",X"09",X"05",X"35",X"32",X"33",
		X"FF",X"82",X"01",X"01",X"16",X"9F",X"AE",X"30",X"19",X"20",X"24",X"34",X"1A",X"21",X"26",X"37",
		X"1B",X"22",X"28",X"FF",X"01",X"01",X"04",X"33",X"9F",X"02",X"00",X"04",X"84",X"9F",X"84",X"01",
		X"04",X"BC",X"9F",X"AD",X"40",X"D1",X"40",X"D1",X"40",X"D1",X"42",X"D1",X"42",X"D1",X"42",X"D1",
		X"39",X"D1",X"39",X"D1",X"39",X"D1",X"39",X"D1",X"3A",X"D1",X"39",X"D1",X"35",X"D1",X"35",X"D1",
		X"35",X"D1",X"35",X"D1",X"34",X"D1",X"32",X"D1",X"30",X"BA",X"D1",X"30",X"D1",X"32",X"D1",X"34",
		X"D1",X"35",X"D1",X"37",X"D1",X"39",X"D1",X"3A",X"D1",X"D2",X"37",X"D1",X"40",X"B4",X"D1",X"40",
		X"D1",X"42",X"D1",X"40",X"D1",X"3A",X"D1",X"39",X"D1",X"37",X"D1",X"35",X"D1",X"D2",X"37",X"D1",
		X"35",X"B4",X"D1",X"FF",X"AE",X"25",X"B4",X"D1",X"29",X"B4",X"D1",X"30",X"B4",X"D1",X"27",X"B4",
		X"D1",X"25",X"B4",X"D1",X"24",X"B4",X"D1",X"22",X"B4",X"D1",X"20",X"B4",X"D1",X"20",X"B4",X"D1",
		X"22",X"B4",X"D1",X"24",X"B4",X"D1",X"20",X"B4",X"D1",X"20",X"D1",X"D2",X"1A",X"D1",X"19",X"D1",
		X"D2",X"17",X"D1",X"15",X"D1",X"D2",X"20",X"D1",X"15",X"B4",X"D1",X"FF",X"AC",X"D4",X"30",X"D5",
		X"30",X"D5",X"30",X"D5",X"30",X"D1",X"D4",X"30",X"D5",X"32",X"D1",X"30",X"D1",X"2A",X"D1",X"29",
		X"D1",X"27",X"D1",X"27",X"D1",X"2B",X"D1",X"32",X"D1",X"34",X"D1",X"35",X"D1",X"37",X"D1",X"39",
		X"D1",X"3A",X"D1",X"40",X"D1",X"D2",X"42",X"D1",X"40",X"B4",X"D1",X"44",X"D1",X"42",X"D1",X"40",
		X"D1",X"3A",X"D1",X"39",X"D1",X"37",X"D1",X"35",X"D1",X"D2",X"30",X"D1",X"35",X"B4",X"D1",X"FF",
		X"D7",X"FF",X"DF",X"5F",X"F7",X"D7",X"FF",X"FF",X"39",X"F7",X"AD",X"5F",X"57",X"57",X"57",X"57",
		X"53",X"57",X"57",X"53",X"57",X"57",X"57",X"57",X"57",X"57",X"4F",X"5F",X"47",X"5F",X"5F",X"47",
		X"47",X"47",X"57",X"47",X"47",X"57",X"47",X"57",X"57",X"47",X"57",X"57",X"57",X"39",X"3F",X"D7",
		X"39",X"3B",X"37",X"36",X"35",X"37",X"36",X"35",X"FF",X"AD",X"55",X"54",X"53",X"52",X"51",X"57",
		X"53",X"57",X"57",X"4B",X"4B",X"57",X"4B",X"4F",X"4B",X"5F",X"47",X"47",X"5F",X"47",X"47",X"47",
		X"47",X"47",X"47",X"57",X"43",X"57",X"57",X"57",X"57",X"57",X"57",X"57",X"57",X"57",X"3B",X"3A",
		X"39",X"3B",X"3A",X"39",X"38",X"37",X"39",X"FF",X"57",X"D7",X"57",X"72",X"A7",X"D7",X"D7",X"57",
		X"78",X"A7",X"E8",X"27",X"5F",X"27",X"B3",X"FF",X"E8",X"21",X"08",X"30",X"B3",X"FF",X"C4",X"01",
		X"01",X"83",X"A0",X"AF",X"33",X"30",X"34",X"31",X"35",X"32",X"36",X"33",X"37",X"34",X"38",X"35",
		X"39",X"36",X"3A",X"37",X"3B",X"FF",X"57",X"DF",X"57",X"A7",X"A7",X"D7",X"57",X"57",X"DE",X"E7",
		X"AD",X"57",X"47",X"47",X"D1",X"47",X"57",X"37",X"D1",X"47",X"47",X"57",X"D1",X"57",X"47",X"D1",
		X"57",X"47",X"D1",X"57",X"47",X"47",X"D1",X"47",X"57",X"37",X"D1",X"47",X"47",X"57",X"D1",X"57",
		X"47",X"D1",X"57",X"47",X"D1",X"57",X"47",X"47",X"D1",X"47",X"57",X"37",X"D1",X"47",X"47",X"57",
		X"D1",X"57",X"47",X"D1",X"57",X"47",X"D1",X"A7",X"E9",X"15",X"15",X"57",X"BF",X"FF",X"AD",X"40",
		X"47",X"44",X"D1",X"44",X"40",X"37",X"D1",X"47",X"44",X"40",X"D1",X"50",X"47",X"D1",X"50",X"47",
		X"D1",X"40",X"47",X"44",X"D1",X"44",X"40",X"37",X"D1",X"47",X"44",X"40",X"D1",X"50",X"47",X"D1",
		X"50",X"47",X"D1",X"40",X"47",X"44",X"D1",X"44",X"40",X"37",X"D1",X"47",X"44",X"40",X"D1",X"50",
		X"47",X"D1",X"50",X"47",X"D1",X"A0",X"E9",X"15",X"15",X"50",X"BF",X"FF",X"42",X"00",X"03",X"26",
		X"A1",X"C4",X"00",X"03",X"3B",X"A2",X"AB",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",
		X"39",X"B2",X"D1",X"3B",X"B2",X"D1",X"39",X"B2",X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"34",
		X"B2",X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"34",X"B2",X"D1",X"32",X"BA",X"D5",X"37",X"B2",
		X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"39",X"B2",X"D1",X"3B",X"B2",X"D1",X"39",X"B2",X"D1",
		X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"44",X"B2",X"D1",X"44",X"B2",X"D1",X"44",X"B2",X"D1",X"44",
		X"B2",X"D1",X"42",X"BA",X"D5",X"3B",X"B2",X"D1",X"3B",X"B2",X"D1",X"3B",X"B2",X"D1",X"3B",X"B2",
		X"D1",X"3B",X"B2",X"D1",X"39",X"B2",X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"32",X"B2",X"D1",
		X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"39",X"B2",X"D1",X"3B",X"BA",X"D5",X"44",X"B6",X"D1",X"44",
		X"B2",X"D1",X"44",X"B2",X"D1",X"42",X"B3",X"37",X"B2",X"D1",X"37",X"B3",X"37",X"B2",X"D1",X"39",
		X"B2",X"D1",X"40",X"B2",X"D1",X"3B",X"B2",X"D1",X"39",X"B2",X"D1",X"37",X"BA",X"D5",X"42",X"B2",
		X"D1",X"42",X"B2",X"D1",X"42",X"B6",X"D1",X"42",X"B2",X"D1",X"42",X"B2",X"D1",X"42",X"B6",X"D1",
		X"44",X"B6",X"D1",X"44",X"B2",X"D1",X"44",X"B3",X"42",X"BA",X"D5",X"44",X"B6",X"D1",X"44",X"B2",
		X"D1",X"44",X"B2",X"D1",X"42",X"B2",X"D1",X"42",X"B2",X"D1",X"42",X"B2",X"D1",X"3B",X"B2",X"D1",
		X"39",X"B2",X"D1",X"39",X"B2",X"D1",X"39",X"B2",X"D1",X"39",X"B2",X"D1",X"42",X"BA",X"D5",X"42",
		X"B2",X"D1",X"42",X"B2",X"D1",X"42",X"B6",X"D1",X"42",X"B2",X"D1",X"42",X"B2",X"D1",X"42",X"B6",
		X"D1",X"44",X"B6",X"D1",X"44",X"B2",X"D1",X"44",X"B3",X"42",X"BA",X"D5",X"44",X"B6",X"D1",X"44",
		X"B2",X"D1",X"44",X"B2",X"D1",X"42",X"B6",X"D1",X"3B",X"B2",X"D1",X"3B",X"B2",X"D1",X"39",X"B6",
		X"D1",X"3B",X"B2",X"D1",X"39",X"B2",X"D1",X"37",X"BA",X"D5",X"FF",X"AA",X"27",X"B2",X"D1",X"3B",
		X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"3B",X"D1",X"42",
		X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"24",
		X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",
		X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",
		X"42",X"D1",X"27",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",
		X"27",X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"24",X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"22",X"B2",
		X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"3B",
		X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"3B",X"D1",X"42",
		X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"24",
		X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",
		X"3B",X"D1",X"42",X"D1",X"27",X"B2",X"D1",X"40",X"D1",X"44",X"D1",X"24",X"B2",X"D1",X"40",X"D1",
		X"44",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",X"22",X"B2",X"D1",X"3B",X"D1",X"42",X"D1",
		X"22",X"B2",X"D1",X"39",X"D1",X"40",X"D1",X"24",X"B2",X"D1",X"25",X"B2",X"D1",X"27",X"B2",X"D1",
		X"22",X"B2",X"D1",X"24",X"B2",X"D1",X"25",X"B2",X"D1",X"27",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",
		X"B2",X"D1",X"2B",X"B2",X"D1",X"27",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",X"B2",X"D1",X"2B",X"B2",
		X"D1",X"34",X"B2",X"D1",X"30",X"B2",X"D1",X"27",X"B2",X"D1",X"34",X"B2",X"D1",X"27",X"B2",X"D1",
		X"2B",X"B2",X"D1",X"32",X"B2",X"D1",X"2B",X"B2",X"D1",X"34",X"B2",X"D1",X"32",X"B2",X"D1",X"30",
		X"B2",X"D1",X"34",X"B2",X"D1",X"32",X"B2",X"D1",X"30",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",X"B2",
		X"D1",X"39",X"B2",X"D1",X"2B",X"B2",X"D1",X"30",X"B2",X"D1",X"31",X"B2",X"D1",X"32",X"B2",X"D1",
		X"22",X"B2",X"D1",X"24",X"B2",X"D1",X"26",X"B2",X"D1",X"27",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",
		X"B2",X"D1",X"2B",X"B2",X"D1",X"27",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",X"B2",X"D1",X"2B",X"B2",
		X"D1",X"34",X"B2",X"D1",X"30",X"B2",X"D1",X"27",X"B2",X"D1",X"34",X"B2",X"D1",X"27",X"B2",X"D1",
		X"2B",X"B2",X"D1",X"32",X"B2",X"D1",X"2B",X"B2",X"D1",X"34",X"B2",X"D1",X"32",X"B2",X"D1",X"30",
		X"B2",X"D1",X"34",X"B2",X"D1",X"32",X"B2",X"D1",X"30",X"B2",X"D1",X"2B",X"B2",X"D1",X"32",X"B2",
		X"D1",X"39",X"B2",X"D1",X"22",X"B2",X"D1",X"24",X"B2",X"D1",X"26",X"B2",X"D1",X"27",X"B2",X"D5",
		X"22",X"B6",X"D1",X"FF",X"C1",X"00",X"02",X"D9",X"A3",X"E8",X"01",X"01",X"C0",X"02",X"BF",X"90",
		X"C1",X"FF",X"81",X"00",X"04",X"E7",X"A3",X"E8",X"10",X"05",X"C0",X"05",X"60",X"90",X"C1",X"D1",
		X"E9",X"10",X"25",X"C0",X"05",X"63",X"BF",X"B8",X"FF",X"C1",X"00",X"03",X"FE",X"A3",X"B2",X"E8",
		X"10",X"02",X"C0",X"10",X"68",X"B9",X"FF",X"02",X"00",X"04",X"11",X"A4",X"84",X"00",X"04",X"1B",
		X"A4",X"E9",X"10",X"20",X"5B",X"56",X"53",X"57",X"BF",X"B6",X"FF",X"E9",X"10",X"20",X"66",X"62",
		X"68",X"61",X"BF",X"B6",X"FF",X"81",X"00",X"03",X"2A",X"A4",X"AD",X"51",X"4A",X"D1",X"51",X"4A",
		X"51",X"4A",X"D1",X"51",X"4A",X"D1",X"51",X"4A",X"51",X"4A",X"D1",X"51",X"4A",X"D1",X"51",X"4A",
		X"51",X"4A",X"D1",X"51",X"4A",X"D1",X"51",X"4A",X"51",X"4A",X"D1",X"51",X"4A",X"D1",X"51",X"4A",
		X"51",X"4A",X"D1",X"51",X"4A",X"D1",X"51",X"4A",X"51",X"4A",X"D1",X"FF",X"C1",X"00",X"03",X"61",
		X"A4",X"AB",X"50",X"54",X"D1",X"50",X"54",X"D1",X"FF",X"02",X"01",X"02",X"73",X"A4",X"84",X"01",
		X"02",X"93",X"A4",X"AD",X"37",X"B2",X"D1",X"36",X"B2",X"D1",X"37",X"B2",X"D1",X"39",X"B2",X"D1",
		X"3B",X"B2",X"D1",X"39",X"B2",X"D1",X"3B",X"B2",X"D1",X"40",X"B2",X"D1",X"42",X"BD",X"D1",X"32",
		X"BD",X"D1",X"FF",X"AD",X"34",X"B2",X"D1",X"33",X"B2",X"D1",X"34",X"B2",X"D1",X"36",X"B2",X"D1",
		X"37",X"B2",X"D1",X"36",X"B2",X"D1",X"37",X"B2",X"D1",X"37",X"B2",X"D1",X"39",X"BD",X"D1",X"29",
		X"BD",X"D1",X"FF",X"01",X"00",X"03",X"BD",X"A4",X"82",X"00",X"03",X"C6",X"A4",X"E9",X"20",X"20",
		X"C0",X"15",X"BF",X"90",X"C1",X"FF",X"E9",X"20",X"20",X"C0",X"15",X"BF",X"90",X"C1",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"A0",X"4D",X"21",X"00",X"4B",X"06",X"02",X"CF",X"3E",X"23",X"06",X"04",X"FF",X"3E",X"10",
		X"CD",X"27",X"A5",X"3A",X"00",X"4B",X"3C",X"FE",X"04",X"38",X"01",X"AF",X"32",X"00",X"4B",X"3E",
		X"0E",X"CD",X"27",X"A5",X"C3",X"09",X"A5",X"F5",X"21",X"5E",X"45",X"3A",X"00",X"4B",X"06",X"0C",
		X"B7",X"28",X"07",X"05",X"3D",X"CD",X"79",X"90",X"18",X"F6",X"F1",X"0E",X"01",X"0D",X"20",X"03",
		X"0E",X"04",X"77",X"05",X"28",X"05",X"CD",X"79",X"90",X"18",X"F2",X"2B",X"06",X"02",X"0D",X"20",
		X"03",X"0E",X"04",X"77",X"05",X"28",X"03",X"2B",X"18",X"F4",X"11",X"E0",X"FF",X"19",X"06",X"0B",
		X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"28",X"06",X"11",X"E0",X"FF",X"19",X"18",X"F1",X"23",
		X"06",X"02",X"0D",X"20",X"03",X"0E",X"04",X"77",X"05",X"C8",X"23",X"18",X"F5",X"FF",X"FF",X"FF",
		X"DD",X"21",X"D4",X"A5",X"CD",X"0A",X"8F",X"DD",X"21",X"F6",X"40",X"FD",X"21",X"F0",X"A5",X"06",
		X"09",X"C5",X"DD",X"E5",X"E1",X"FD",X"7E",X"00",X"FD",X"5E",X"01",X"01",X"02",X"02",X"CD",X"5C",
		X"90",X"DD",X"E5",X"E1",X"11",X"40",X"00",X"19",X"3E",X"3A",X"1E",X"00",X"01",X"04",X"01",X"CD",
		X"4A",X"90",X"DD",X"E5",X"FD",X"6E",X"02",X"FD",X"66",X"03",X"E5",X"DD",X"E1",X"CD",X"0A",X"8F",
		X"3E",X"23",X"06",X"08",X"FF",X"11",X"04",X"00",X"FD",X"19",X"DD",X"E1",X"DD",X"2B",X"DD",X"2B",
		X"C1",X"10",X"BE",X"C9",X"00",X"05",X"BC",X"41",X"01",X"02",X"44",X"14",X"52",X"03",X"45",X"04",
		X"41",X"05",X"4D",X"07",X"9A",X"41",X"00",X"05",X"53",X"48",X"4F",X"50",X"50",X"45",X"52",X"00",
		X"B8",X"0D",X"14",X"A6",X"B8",X"0E",X"26",X"A6",X"B8",X"0F",X"38",X"A6",X"B8",X"10",X"4A",X"A6",
		X"C0",X"0D",X"5C",X"A6",X"C4",X"0E",X"6A",X"A6",X"C8",X"0F",X"78",X"A6",X"CC",X"10",X"86",X"A6",
		X"01",X"0A",X"94",X"A6",X"04",X"0B",X"D6",X"41",X"00",X"02",X"4D",X"49",X"53",X"54",X"45",X"52",
		X"59",X"20",X"50",X"54",X"53",X"00",X"04",X"0B",X"D4",X"41",X"00",X"03",X"4D",X"49",X"53",X"54",
		X"45",X"52",X"59",X"20",X"50",X"54",X"53",X"00",X"04",X"0B",X"D2",X"41",X"00",X"04",X"4D",X"49",
		X"53",X"54",X"45",X"52",X"59",X"20",X"50",X"54",X"53",X"00",X"04",X"0B",X"D0",X"41",X"00",X"05",
		X"4D",X"49",X"53",X"54",X"45",X"52",X"59",X"20",X"50",X"54",X"53",X"00",X"04",X"07",X"CE",X"41",
		X"00",X"02",X"35",X"30",X"30",X"20",X"50",X"54",X"53",X"00",X"04",X"07",X"CC",X"41",X"00",X"03",
		X"32",X"35",X"30",X"20",X"50",X"54",X"53",X"00",X"04",X"07",X"CA",X"41",X"00",X"04",X"31",X"30",
		X"30",X"20",X"50",X"54",X"53",X"00",X"04",X"07",X"C8",X"41",X"00",X"05",X"20",X"35",X"30",X"20",
		X"50",X"54",X"53",X"00",X"04",X"04",X"C6",X"41",X"00",X"04",X"42",X"4F",X"4D",X"42",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"C0",X"4F",X"AF",X"32",X"C0",X"50",X"1E",X"00",X"21",X"00",X"40",X"01",X"00",X"10",X"73",
		X"23",X"0D",X"20",X"FB",X"AF",X"32",X"C0",X"50",X"10",X"F5",X"21",X"00",X"40",X"01",X"00",X"10",
		X"7E",X"BB",X"20",X"15",X"23",X"0D",X"20",X"F8",X"AF",X"32",X"C0",X"50",X"10",X"F2",X"3E",X"11",
		X"83",X"5F",X"E6",X"0F",X"20",X"D3",X"C3",X"60",X"A7",X"AF",X"32",X"C0",X"50",X"DD",X"21",X"78",
		X"A7",X"7C",X"FE",X"48",X"38",X"04",X"DD",X"21",X"8A",X"A7",X"CD",X"0A",X"8F",X"AF",X"32",X"C0",
		X"50",X"01",X"00",X"00",X"0D",X"20",X"FD",X"AF",X"32",X"C0",X"50",X"10",X"F7",X"C3",X"03",X"A7",
		X"21",X"02",X"48",X"CB",X"66",X"CB",X"E6",X"EF",X"CD",X"07",X"AC",X"DD",X"21",X"9C",X"A7",X"CD",
		X"0A",X"8F",X"CD",X"11",X"AC",X"C3",X"AF",X"A7",X"00",X"0B",X"4F",X"41",X"00",X"00",X"52",X"41",
		X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"3B",X"31",X"00",X"00",X"0B",X"4F",X"41",X"00",X"00",
		X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"3B",X"32",X"00",X"00",X"0C",X"4F",X"41",
		X"00",X"05",X"52",X"41",X"4D",X"20",X"43",X"48",X"45",X"43",X"4B",X"20",X"4F",X"4B",X"00",X"CD",
		X"07",X"AC",X"DD",X"21",X"1F",X"A8",X"CD",X"0A",X"8F",X"DD",X"21",X"95",X"41",X"21",X"00",X"00",
		X"11",X"2F",X"A8",X"AF",X"01",X"00",X"10",X"86",X"23",X"0D",X"20",X"FB",X"10",X"F9",X"47",X"1A",
		X"B8",X"CD",X"ED",X"A7",X"DD",X"2B",X"DD",X"2B",X"13",X"7C",X"FE",X"B0",X"28",X"09",X"FE",X"40",
		X"20",X"E1",X"21",X"00",X"80",X"18",X"DC",X"CD",X"11",X"AC",X"C3",X"47",X"A8",X"06",X"08",X"E5",
		X"D5",X"DD",X"E5",X"E1",X"11",X"37",X"A8",X"28",X"03",X"11",X"3F",X"A8",X"1A",X"77",X"13",X"CD",
		X"79",X"90",X"10",X"F8",X"E1",X"E5",X"01",X"2F",X"A8",X"B7",X"ED",X"42",X"7D",X"3C",X"F6",X"30",
		X"DD",X"E5",X"11",X"80",X"00",X"DD",X"19",X"DD",X"77",X"00",X"DD",X"E1",X"D1",X"E1",X"C9",X"00",
		X"09",X"9A",X"41",X"00",X"17",X"52",X"4F",X"4D",X"20",X"43",X"48",X"45",X"43",X"4B",X"00",X"FE",
		X"74",X"94",X"D1",X"2F",X"7D",X"00",X"42",X"52",X"4F",X"4D",X"3B",X"20",X"20",X"4F",X"4B",X"52",
		X"4F",X"4D",X"3B",X"20",X"42",X"41",X"44",X"CD",X"07",X"AC",X"DD",X"21",X"49",X"A9",X"CD",X"0A",
		X"8F",X"DD",X"21",X"04",X"AA",X"CD",X"0A",X"8F",X"3A",X"00",X"50",X"2F",X"E6",X"BF",X"21",X"DC",
		X"44",X"CD",X"F4",X"A8",X"3A",X"40",X"50",X"2F",X"E6",X"7F",X"FE",X"60",X"CA",X"0E",X"A9",X"21",
		X"3C",X"46",X"CD",X"F4",X"A8",X"3A",X"80",X"50",X"2F",X"21",X"0F",X"45",X"06",X"08",X"1E",X"00",
		X"CB",X"3F",X"30",X"02",X"1E",X"04",X"73",X"CD",X"79",X"90",X"CD",X"79",X"90",X"10",X"EF",X"3A",
		X"80",X"50",X"2F",X"CB",X"47",X"DD",X"21",X"DA",X"AB",X"20",X"04",X"DD",X"21",X"E9",X"AB",X"F5",
		X"CD",X"0A",X"8F",X"F1",X"F5",X"E6",X"02",X"CB",X"3F",X"32",X"03",X"50",X"F1",X"F5",X"E6",X"0C",
		X"CB",X"3F",X"CB",X"3F",X"21",X"76",X"AA",X"CD",X"1D",X"94",X"D5",X"DD",X"E1",X"CD",X"0A",X"8F",
		X"F1",X"F5",X"E6",X"30",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"C6",X"33",X"21",X"65",
		X"42",X"77",X"CB",X"D4",X"36",X"14",X"F1",X"E6",X"C0",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"76",X"AB",X"CD",X"1D",X"94",X"D5",X"DD",X"E1",X"CD",X"0A",
		X"8F",X"C3",X"58",X"A8",X"06",X"08",X"E5",X"C5",X"1E",X"00",X"CB",X"3F",X"30",X"02",X"1E",X"04",
		X"06",X"09",X"73",X"CD",X"79",X"90",X"10",X"FA",X"C1",X"E1",X"2B",X"10",X"E9",X"C9",X"21",X"00",
		X"40",X"1E",X"16",X"3E",X"00",X"01",X"20",X"20",X"CD",X"4A",X"90",X"3E",X"01",X"32",X"02",X"50",
		X"32",X"01",X"50",X"3A",X"00",X"50",X"2F",X"E6",X"0F",X"28",X"F8",X"11",X"00",X"00",X"FE",X"01",
		X"28",X"11",X"11",X"01",X"00",X"FE",X"02",X"28",X"0A",X"11",X"00",X"01",X"FE",X"04",X"28",X"03",
		X"11",X"01",X"01",X"ED",X"53",X"05",X"50",X"18",X"DA",X"00",X"0E",X"3E",X"41",X"00",X"17",X"43",
		X"4F",X"4E",X"54",X"52",X"4F",X"4C",X"45",X"52",X"20",X"54",X"45",X"53",X"54",X"11",X"DC",X"40",
		X"00",X"00",X"50",X"31",X"3A",X"3A",X"55",X"50",X"20",X"20",X"20",X"20",X"20",X"50",X"32",X"3A",
		X"3A",X"55",X"50",X"13",X"DB",X"40",X"00",X"00",X"50",X"31",X"3A",X"3A",X"4C",X"45",X"46",X"54",
		X"20",X"20",X"20",X"50",X"32",X"3A",X"3A",X"4C",X"45",X"46",X"54",X"14",X"DA",X"40",X"00",X"00",
		X"50",X"31",X"3A",X"3A",X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"50",X"32",X"3A",X"3A",X"52",
		X"49",X"47",X"48",X"54",X"13",X"D9",X"40",X"00",X"00",X"50",X"31",X"3A",X"3A",X"44",X"4F",X"57",
		X"4E",X"20",X"20",X"20",X"50",X"32",X"3A",X"3A",X"44",X"4F",X"57",X"4E",X"13",X"D8",X"40",X"00",
		X"00",X"50",X"31",X"3A",X"3A",X"50",X"55",X"53",X"48",X"20",X"20",X"20",X"50",X"32",X"3A",X"3A",
		X"50",X"55",X"53",X"48",X"11",X"17",X"41",X"00",X"00",X"43",X"4F",X"49",X"4E",X"20",X"20",X"20",
		X"20",X"20",X"31",X"50",X"3A",X"53",X"54",X"41",X"52",X"54",X"08",X"36",X"42",X"00",X"00",X"32",
		X"50",X"3A",X"53",X"54",X"41",X"52",X"54",X"07",X"F5",X"40",X"00",X"00",X"53",X"45",X"52",X"56",
		X"49",X"43",X"45",X"00",X"00",X"0B",X"71",X"41",X"00",X"17",X"44",X"49",X"50",X"3B",X"53",X"57",
		X"20",X"54",X"45",X"53",X"54",X"0F",X"0F",X"41",X"00",X"00",X"31",X"20",X"32",X"20",X"33",X"20",
		X"34",X"20",X"35",X"20",X"36",X"20",X"37",X"20",X"38",X"0E",X"AC",X"40",X"00",X"00",X"47",X"41",
		X"4D",X"45",X"20",X"53",X"54",X"59",X"4C",X"45",X"3A",X"3A",X"3A",X"3A",X"0E",X"AA",X"40",X"00",
		X"00",X"42",X"4F",X"4E",X"55",X"53",X"20",X"4C",X"49",X"56",X"45",X"53",X"3A",X"3A",X"3A",X"0E",
		X"A5",X"40",X"00",X"00",X"43",X"48",X"41",X"52",X"4C",X"45",X"59",X"20",X"4F",X"57",X"4E",X"3A",
		X"3A",X"3A",X"0E",X"A3",X"40",X"00",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"3A",X"3A",X"3A",
		X"3A",X"3A",X"3A",X"3A",X"3A",X"00",X"7E",X"AA",X"BC",X"AA",X"FA",X"AA",X"38",X"AB",X"00",X"0A",
		X"6A",X"42",X"00",X"04",X"4E",X"4F",X"20",X"42",X"4F",X"4E",X"55",X"53",X"20",X"20",X"0A",X"69",
		X"42",X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"0A",X"68",X"42",
		X"00",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"0A",X"67",X"42",X"00",
		X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"00",X"0A",X"6A",X"42",
		X"00",X"05",X"31",X"53",X"54",X"20",X"20",X"33",X"30",X"30",X"30",X"30",X"0A",X"69",X"42",X"00",
		X"04",X"32",X"4E",X"44",X"20",X"20",X"36",X"30",X"30",X"30",X"30",X"0A",X"68",X"42",X"00",X"17",
		X"33",X"52",X"44",X"20",X"31",X"35",X"30",X"30",X"30",X"30",X"0A",X"67",X"42",X"00",X"02",X"34",
		X"54",X"48",X"20",X"32",X"35",X"30",X"30",X"30",X"30",X"00",X"00",X"0A",X"6A",X"42",X"00",X"05",
		X"31",X"53",X"54",X"20",X"20",X"35",X"30",X"30",X"30",X"30",X"0A",X"69",X"42",X"00",X"04",X"32",
		X"4E",X"44",X"20",X"31",X"30",X"30",X"30",X"30",X"30",X"0A",X"68",X"42",X"00",X"17",X"33",X"52",
		X"44",X"20",X"32",X"30",X"30",X"30",X"30",X"30",X"0A",X"67",X"42",X"00",X"02",X"34",X"54",X"48",
		X"20",X"35",X"30",X"30",X"30",X"30",X"30",X"00",X"00",X"0A",X"6A",X"42",X"00",X"05",X"31",X"53",
		X"54",X"20",X"20",X"37",X"30",X"30",X"30",X"30",X"0A",X"69",X"42",X"00",X"04",X"32",X"4E",X"44",
		X"20",X"31",X"35",X"30",X"30",X"30",X"30",X"0A",X"68",X"42",X"00",X"17",X"33",X"52",X"44",X"20",
		X"33",X"30",X"30",X"30",X"30",X"30",X"0A",X"67",X"42",X"00",X"02",X"34",X"54",X"48",X"20",X"37",
		X"30",X"30",X"30",X"30",X"30",X"00",X"7E",X"AB",X"95",X"AB",X"AC",X"AB",X"C3",X"AB",X"00",X"10",
		X"C3",X"41",X"00",X"05",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"31",X"20",X"43",X"52",X"45",
		X"44",X"49",X"54",X"20",X"00",X"00",X"10",X"C3",X"41",X"00",X"05",X"31",X"20",X"43",X"4F",X"49",
		X"4E",X"20",X"32",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"20",X"00",X"00",X"10",X"C3",X"41",
		X"00",X"05",X"31",X"20",X"43",X"4F",X"49",X"4E",X"20",X"33",X"20",X"43",X"52",X"45",X"44",X"49",
		X"54",X"20",X"00",X"00",X"10",X"C3",X"41",X"00",X"05",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",
		X"20",X"31",X"20",X"43",X"52",X"45",X"44",X"49",X"54",X"00",X"00",X"08",X"6C",X"42",X"00",X"04",
		X"54",X"41",X"42",X"4C",X"45",X"20",X"20",X"20",X"00",X"00",X"08",X"6C",X"42",X"00",X"04",X"55",
		X"50",X"20",X"52",X"49",X"47",X"48",X"54",X"00",X"00",X"08",X"6A",X"42",X"00",X"04",X"4E",X"4F",
		X"20",X"42",X"4F",X"4E",X"55",X"53",X"00",X"21",X"00",X"40",X"01",X"00",X"08",X"CD",X"00",X"8F",
		X"C9",X"3E",X"05",X"01",X"FF",X"FF",X"0D",X"20",X"FD",X"05",X"20",X"FA",X"3D",X"20",X"F4",X"C9",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"31",X"20",X"4E",X"21",X"A0",X"4A",X"06",X"1E",X"CF",X"3E",X"23",X"06",X"01",X"FF",X"FD",X"21",
		X"A0",X"4A",X"06",X"03",X"C5",X"FD",X"7E",X"00",X"B7",X"C4",X"26",X"AD",X"01",X"0A",X"00",X"FD",
		X"09",X"C1",X"10",X"F0",X"18",X"E3",X"FE",X"01",X"C2",X"DB",X"AD",X"FD",X"35",X"05",X"C2",X"50",
		X"AD",X"FD",X"34",X"00",X"FD",X"36",X"06",X"00",X"FD",X"36",X"07",X"00",X"FD",X"66",X"01",X"FD",
		X"6E",X"02",X"CD",X"1E",X"92",X"01",X"02",X"02",X"3E",X"09",X"1E",X"0B",X"CD",X"5C",X"90",X"C9",
		X"FD",X"7E",X"07",X"CB",X"BF",X"B7",X"28",X"06",X"FD",X"35",X"07",X"C3",X"A3",X"AD",X"3E",X"02",
		X"FD",X"B6",X"07",X"FD",X"77",X"07",X"FD",X"66",X"03",X"FD",X"6E",X"04",X"CD",X"1E",X"92",X"1E",
		X"0D",X"FD",X"CB",X"07",X"7E",X"FD",X"CB",X"07",X"FE",X"28",X"06",X"FD",X"CB",X"07",X"BE",X"1E",
		X"10",X"01",X"05",X"05",X"C5",X"E5",X"C5",X"E5",X"3E",X"88",X"01",X"02",X"02",X"CD",X"5C",X"90",
		X"E1",X"23",X"23",X"C1",X"10",X"F0",X"E1",X"01",X"40",X"00",X"09",X"C1",X"0D",X"C2",X"84",X"AD",
		X"C3",X"BF",X"AD",X"FD",X"7E",X"06",X"CB",X"BF",X"B7",X"28",X"04",X"FD",X"35",X"06",X"C9",X"3E",
		X"04",X"FD",X"B6",X"06",X"CB",X"7F",X"CB",X"FF",X"28",X"02",X"CB",X"BF",X"FD",X"77",X"06",X"FD",
		X"66",X"01",X"FD",X"6E",X"02",X"CD",X"1E",X"92",X"3E",X"01",X"FD",X"CB",X"06",X"7E",X"28",X"02",
		X"3E",X"05",X"01",X"02",X"02",X"1E",X"0A",X"CD",X"5C",X"90",X"C9",X"3A",X"02",X"48",X"CB",X"77",
		X"CB",X"F7",X"20",X"0C",X"32",X"02",X"48",X"CB",X"6F",X"20",X"05",X"3E",X"1F",X"CD",X"40",X"03",
		X"FD",X"7E",X"06",X"B7",X"28",X"06",X"FD",X"35",X"06",X"C3",X"1A",X"AE",X"FD",X"36",X"06",X"03",
		X"FD",X"66",X"01",X"FD",X"6E",X"02",X"CD",X"1E",X"92",X"7E",X"FE",X"11",X"20",X"02",X"3E",X"05",
		X"C6",X"04",X"1E",X"0B",X"01",X"02",X"02",X"CD",X"5C",X"90",X"FD",X"7E",X"07",X"B7",X"28",X"04",
		X"FD",X"35",X"07",X"C9",X"FD",X"36",X"07",X"03",X"FD",X"66",X"01",X"FD",X"6E",X"02",X"CD",X"1E",
		X"92",X"E5",X"E5",X"FD",X"7E",X"08",X"3D",X"CB",X"7F",X"28",X"02",X"3E",X"03",X"CD",X"56",X"AF",
		X"E1",X"19",X"3E",X"05",X"CD",X"BC",X"AF",X"FD",X"7E",X"08",X"CD",X"56",X"AF",X"E1",X"19",X"3E",
		X"02",X"CD",X"BC",X"AF",X"FD",X"7E",X"08",X"3C",X"FD",X"77",X"08",X"FE",X"04",X"D8",X"FD",X"36",
		X"08",X"00",X"FD",X"34",X"09",X"3E",X"04",X"FD",X"BE",X"09",X"C0",X"FD",X"E5",X"FD",X"66",X"01",
		X"FD",X"6E",X"02",X"CD",X"AC",X"91",X"36",X"20",X"FD",X"66",X"03",X"FD",X"6E",X"04",X"E5",X"CD",
		X"AC",X"91",X"E5",X"FD",X"E1",X"E1",X"CD",X"1E",X"92",X"E5",X"DD",X"E1",X"01",X"05",X"05",X"C5",
		X"FD",X"E5",X"DD",X"E5",X"C5",X"DD",X"E5",X"E1",X"CD",X"83",X"26",X"30",X"0C",X"3E",X"88",X"1E",
		X"03",X"01",X"02",X"02",X"CD",X"5C",X"90",X"18",X"24",X"FD",X"CB",X"00",X"9E",X"21",X"0C",X"AF",
		X"FD",X"7E",X"00",X"CB",X"7F",X"28",X"03",X"21",X"16",X"AF",X"E6",X"70",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"CB",X"3F",X"CD",X"1D",X"94",X"EB",X"11",X"CD",X"AE",X"D5",X"E9",X"FD",X"23",X"DD",
		X"23",X"DD",X"23",X"C1",X"10",X"BE",X"DD",X"E1",X"11",X"40",X"00",X"DD",X"19",X"FD",X"E1",X"11",
		X"0C",X"00",X"FD",X"19",X"C1",X"0D",X"20",X"A7",X"FD",X"E1",X"FD",X"E5",X"E1",X"06",X"0A",X"CF",
		X"FD",X"E5",X"FD",X"21",X"A0",X"4A",X"06",X"03",X"FD",X"7E",X"00",X"B7",X"20",X"0B",X"FD",X"23",
		X"10",X"F6",X"21",X"02",X"48",X"CB",X"76",X"CB",X"B6",X"FD",X"E1",X"C9",X"20",X"AF",X"20",X"AF",
		X"34",X"AF",X"B6",X"2D",X"27",X"AF",X"44",X"AF",X"44",X"AF",X"34",X"AF",X"44",X"AF",X"34",X"AF",
		X"3A",X"01",X"48",X"CB",X"57",X"20",X"13",X"DD",X"E5",X"E1",X"AF",X"1E",X"16",X"01",X"02",X"02",
		X"CD",X"4A",X"90",X"C9",X"1E",X"14",X"3E",X"88",X"18",X"12",X"FD",X"7E",X"00",X"E6",X"07",X"CD",
		X"76",X"95",X"18",X"08",X"FD",X"7E",X"00",X"E6",X"07",X"CD",X"87",X"95",X"DD",X"E5",X"E1",X"01",
		X"02",X"02",X"CD",X"5C",X"90",X"C9",X"21",X"62",X"AF",X"CD",X"0B",X"94",X"46",X"23",X"5E",X"23",
		X"56",X"C9",X"04",X"DF",X"FF",X"06",X"BE",X"FF",X"08",X"9D",X"FF",X"0A",X"7C",X"FF",X"3E",X"18",
		X"CD",X"40",X"03",X"FD",X"21",X"A0",X"4A",X"06",X"03",X"C5",X"FD",X"7E",X"00",X"B7",X"20",X"33",
		X"FD",X"34",X"00",X"FD",X"74",X"01",X"FD",X"75",X"02",X"3E",X"40",X"FD",X"77",X"05",X"01",X"E0",
		X"20",X"CD",X"A5",X"91",X"FD",X"74",X"03",X"FD",X"75",X"04",X"CD",X"AC",X"91",X"01",X"05",X"05",
		X"C5",X"E5",X"CB",X"DE",X"23",X"10",X"FB",X"E1",X"01",X"0C",X"00",X"09",X"C1",X"0D",X"C2",X"A0",
		X"AF",X"C1",X"C9",X"01",X"0A",X"00",X"FD",X"09",X"C1",X"10",X"BE",X"C9",X"C5",X"CD",X"E6",X"AF",
		X"23",X"10",X"FA",X"2B",X"C1",X"C5",X"11",X"20",X"00",X"CD",X"E6",X"AF",X"19",X"10",X"FA",X"C1",
		X"C5",X"B7",X"ED",X"52",X"CD",X"E6",X"AF",X"2B",X"10",X"FA",X"C1",X"23",X"11",X"E0",X"FF",X"CD",
		X"E6",X"AF",X"19",X"10",X"FA",X"C9",X"36",X"1F",X"CB",X"D4",X"77",X"CB",X"94",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
