library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"F0",X"87",X"3C",X"4B",X"0F",X"0F",X"00",X"70",X"70",X"70",X"70",X"61",X"61",X"61",
		X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"F0",X"F0",X"78",X"3C",X"1E",X"1E",X"1E",
		X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"F0",X"00",X"61",X"61",X"61",X"70",X"70",X"70",X"70",X"00",
		X"68",X"2C",X"A4",X"E4",X"E8",X"E0",X"E0",X"00",X"0F",X"1E",X"1E",X"3C",X"78",X"F2",X"F0",X"00",
		X"00",X"F0",X"F0",X"87",X"3C",X"4B",X"0F",X"0F",X"00",X"70",X"70",X"70",X"70",X"61",X"61",X"61",
		X"00",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"F0",X"F0",X"78",X"3C",X"1E",X"1E",X"1E",
		X"0F",X"0F",X"0F",X"0F",X"87",X"F0",X"F0",X"00",X"61",X"61",X"61",X"70",X"70",X"70",X"70",X"00",
		X"68",X"2C",X"A4",X"E4",X"E0",X"E4",X"E0",X"00",X"0F",X"1E",X"1E",X"3C",X"79",X"F0",X"F0",X"00",
		X"00",X"20",X"11",X"00",X"99",X"CB",X"BC",X"71",X"00",X"00",X"00",X"11",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"44",X"88",X"00",X"00",X"00",X"00",X"00",X"88",X"58",X"87",X"79",X"2C",
		X"BC",X"0F",X"5B",X"20",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"22",X"00",X"10",X"00",X"00",
		X"00",X"80",X"44",X"00",X"00",X"00",X"00",X"00",X"E9",X"96",X"E2",X"0C",X"80",X"40",X"00",X"00",
		X"00",X"01",X"32",X"91",X"4B",X"CC",X"ED",X"4C",X"00",X"00",X"12",X"10",X"33",X"01",X"00",X"01",
		X"00",X"00",X"A8",X"4C",X"08",X"00",X"00",X"00",X"00",X"00",X"80",X"0D",X"69",X"F2",X"CF",X"8E",
		X"C1",X"DC",X"AD",X"0F",X"B2",X"01",X"00",X"00",X"01",X"12",X"11",X"32",X"01",X"50",X"00",X"00",
		X"00",X"08",X"48",X"08",X"88",X"04",X"00",X"00",X"52",X"FC",X"67",X"96",X"3A",X"11",X"00",X"00",
		X"11",X"20",X"C0",X"A6",X"6E",X"7B",X"2C",X"9C",X"80",X"40",X"02",X"21",X"10",X"25",X"21",X"30",
		X"20",X"60",X"0E",X"C0",X"40",X"00",X"00",X"10",X"00",X"00",X"14",X"C3",X"A1",X"67",X"62",X"21",
		X"0F",X"85",X"5E",X"9D",X"0E",X"C0",X"00",X"80",X"10",X"21",X"71",X"53",X"30",X"81",X"32",X"00",
		X"28",X"48",X"C0",X"08",X"40",X"80",X"20",X"10",X"D2",X"07",X"E7",X"ED",X"43",X"C2",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"00",X"00",X"44",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"11",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"FF",
		X"00",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"48",X"00",X"00",X"00",X"08",X"0E",X"0F",X"6F",X"8F",
		X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"60",X"60",X"00",X"00",X"00",
		X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",X"FF",X"88",X"CC",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"EE",X"CC",X"88",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",X"8F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"60",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"68",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"6F",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"60",X"60",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"48",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"8F",X"6F",X"0F",X"0E",X"08",X"00",X"00",X"00",
		X"00",X"C3",X"C3",X"F0",X"F0",X"F2",X"F6",X"FE",X"00",X"04",X"12",X"16",X"16",X"34",X"70",X"30",
		X"00",X"80",X"C0",X"C0",X"C0",X"0E",X"48",X"E0",X"00",X"78",X"F0",X"F0",X"F6",X"F7",X"2F",X"BD",
		X"FE",X"F6",X"F2",X"F0",X"F0",X"C3",X"C3",X"00",X"30",X"70",X"34",X"16",X"16",X"12",X"04",X"00",
		X"E0",X"48",X"0E",X"C0",X"C0",X"C0",X"80",X"00",X"BD",X"2F",X"F7",X"F6",X"F0",X"F0",X"78",X"00",
		X"44",X"5F",X"5F",X"D7",X"5F",X"D7",X"44",X"00",X"0C",X"2D",X"3C",X"78",X"3C",X"38",X"10",X"00",
		X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"C3",X"CB",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"3C",X"3D",
		X"CB",X"C3",X"0F",X"0F",X"0F",X"0F",X"C3",X"CB",X"3D",X"3C",X"0F",X"0F",X"0F",X"0F",X"3C",X"3D",
		X"00",X"CC",X"EE",X"11",X"11",X"33",X"EE",X"CC",X"00",X"11",X"33",X"66",X"44",X"44",X"33",X"11",
		X"00",X"00",X"00",X"22",X"FF",X"FF",X"00",X"00",X"00",X"00",X"44",X"44",X"77",X"77",X"44",X"44",
		X"00",X"22",X"33",X"99",X"99",X"DD",X"FF",X"66",X"00",X"66",X"77",X"77",X"55",X"55",X"44",X"44",
		X"00",X"00",X"11",X"99",X"DD",X"FF",X"BB",X"11",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"88",X"CC",X"66",X"33",X"FF",X"FF",X"00",X"00",X"11",X"11",X"11",X"11",X"77",X"77",X"11",
		X"00",X"77",X"77",X"55",X"55",X"55",X"DD",X"88",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"CC",X"EE",X"BB",X"99",X"99",X"99",X"00",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"33",X"33",X"11",X"99",X"DD",X"77",X"33",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"00",
		X"00",X"66",X"FF",X"DD",X"99",X"99",X"66",X"00",X"00",X"33",X"44",X"44",X"55",X"55",X"77",X"33",
		X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"EE",X"00",X"00",X"44",X"44",X"44",X"66",X"33",X"11",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"00",
		X"00",X"00",X"88",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CB",X"C3",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"3D",X"3C",X"0F",X"0F",X"0F",X"0F",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"33",X"11",X"99",X"DD",X"99",X"BB",X"EE",X"77",X"CC",X"88",X"99",X"BB",X"99",X"DD",X"77",
		X"00",X"CC",X"EE",X"33",X"11",X"33",X"EE",X"CC",X"00",X"77",X"77",X"11",X"11",X"11",X"77",X"77",
		X"00",X"FF",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",X"77",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"CC",X"EE",X"33",X"11",X"11",X"33",X"22",X"00",X"11",X"33",X"66",X"44",X"44",X"66",X"22",
		X"00",X"FF",X"FF",X"11",X"11",X"33",X"EE",X"CC",X"00",X"77",X"77",X"44",X"44",X"66",X"33",X"11",
		X"00",X"00",X"FF",X"FF",X"99",X"99",X"99",X"11",X"00",X"00",X"77",X"77",X"44",X"44",X"44",X"44",
		X"00",X"FF",X"FF",X"99",X"99",X"99",X"99",X"11",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CC",X"EE",X"33",X"11",X"99",X"99",X"99",X"00",X"11",X"33",X"66",X"44",X"44",X"77",X"77",
		X"00",X"FF",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",X"77",X"77",X"00",X"00",X"00",X"77",X"77",
		X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"44",X"44",X"77",X"77",X"44",X"44",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"22",X"66",X"44",X"44",X"66",X"77",X"33",
		X"00",X"FF",X"FF",X"88",X"CC",X"66",X"33",X"11",X"00",X"77",X"77",X"11",X"33",X"77",X"66",X"44",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"44",X"44",X"44",X"44",
		X"00",X"FF",X"FF",X"EE",X"CC",X"EE",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"00",X"77",X"77",
		X"00",X"FF",X"FF",X"EE",X"CC",X"88",X"FF",X"FF",X"00",X"77",X"77",X"00",X"11",X"33",X"77",X"77",
		X"00",X"EE",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"EE",X"00",X"77",X"77",X"11",X"11",X"11",X"11",X"00",
		X"F0",X"F0",X"78",X"3C",X"3C",X"78",X"F0",X"F0",X"F0",X"F0",X"E1",X"C3",X"C3",X"E1",X"F0",X"F0",
		X"00",X"FF",X"FF",X"11",X"11",X"99",X"FF",X"EE",X"00",X"77",X"77",X"11",X"33",X"77",X"66",X"44",
		X"00",X"66",X"FF",X"99",X"99",X"BB",X"AA",X"00",X"00",X"22",X"66",X"44",X"44",X"44",X"77",X"33",
		X"00",X"00",X"11",X"11",X"FF",X"FF",X"11",X"11",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",X"33",X"77",X"44",X"44",X"44",X"77",X"33",
		X"00",X"FF",X"FF",X"88",X"00",X"88",X"FF",X"FF",X"00",X"00",X"11",X"33",X"77",X"33",X"11",X"00",
		X"00",X"FF",X"FF",X"88",X"CC",X"88",X"FF",X"FF",X"00",X"11",X"77",X"33",X"11",X"33",X"77",X"11",
		X"00",X"33",X"77",X"EE",X"CC",X"EE",X"77",X"33",X"00",X"66",X"77",X"33",X"11",X"33",X"77",X"66",
		X"00",X"00",X"33",X"FF",X"88",X"88",X"FF",X"33",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"00",
		X"00",X"11",X"11",X"99",X"DD",X"FF",X"77",X"33",X"00",X"66",X"77",X"77",X"55",X"44",X"44",X"44",
		X"00",X"00",X"88",X"CC",X"66",X"33",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"66",X"00",X"00",
		X"FA",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"33",X"66",X"CC",X"88",X"00",X"00",X"00",X"00",X"66",X"33",X"11",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"FF",X"FF",X"CF",X"0F",X"0F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"EF",X"EF",X"CF",X"CF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"0F",X"2F",X"4F",X"5F",
		X"0F",X"0F",X"4F",X"3F",X"0F",X"CF",X"FF",X"FF",X"CF",X"CF",X"EF",X"EF",X"FF",X"FF",X"FF",X"FF",
		X"F7",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"5E",X"1F",X"0F",X"0F",X"1F",X"3F",X"FF",X"FF",
		X"00",X"00",X"11",X"11",X"75",X"FF",X"F7",X"FE",X"00",X"00",X"00",X"32",X"33",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"80",X"88",X"EC",X"E6",X"FA",X"FF",
		X"FF",X"FD",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"EF",X"F7",X"EE",X"FB",X"CC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"78",X"A5",X"4B",X"B4",X"96",X"00",X"00",X"00",X"00",X"10",X"12",X"21",X"03",
		X"00",X"00",X"00",X"00",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"00",X"80",X"C0",X"84",X"48",
		X"5A",X"96",X"4B",X"A5",X"96",X"0F",X"00",X"00",X"12",X"12",X"03",X"12",X"01",X"00",X"00",X"00",
		X"08",X"08",X"0C",X"04",X"04",X"00",X"00",X"00",X"85",X"0E",X"84",X"0C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"02",X"74",X"74",X"74",X"F4",X"F4",X"00",X"00",X"00",X"02",X"32",X"32",X"32",X"32",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"F2",X"F1",X"F8",X"FC",X"77",X"00",X"00",X"00",X"32",X"33",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"08",X"08",X"08",X"00",X"00",X"00",X"C0",X"E0",X"F8",X"E1",X"CA",X"00",X"00",X"00",
		X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",
		X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"10",X"31",X"73",X"F7",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"10",X"31",X"73",X"F7",
		X"00",X"00",X"00",X"00",X"80",X"C8",X"EC",X"FE",X"80",X"C8",X"EC",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",
		X"FE",X"EC",X"C8",X"80",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FE",X"EC",X"C8",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"F7",X"73",X"31",X"10",X"F7",X"73",X"31",X"10",X"00",X"00",X"00",X"00",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FA",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F5",
		X"F5",X"FE",X"EC",X"C8",X"80",X"00",X"00",X"00",X"F5",X"FF",X"FF",X"FF",X"FF",X"FE",X"EC",X"C8",
		X"FE",X"FF",X"FE",X"FF",X"FE",X"FF",X"FE",X"F5",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F5",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",
		X"FA",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FA",X"F7",X"FF",X"F7",X"FF",X"F7",X"FF",X"F7",
		X"00",X"00",X"00",X"00",X"80",X"E6",X"E6",X"E6",X"C0",X"C0",X"E0",X"70",X"30",X"10",X"F0",X"30",
		X"EE",X"11",X"11",X"22",X"22",X"11",X"11",X"EE",X"11",X"C3",X"C3",X"E7",X"E7",X"C3",X"C3",X"11",
		X"CC",X"22",X"11",X"11",X"11",X"11",X"66",X"88",X"E0",X"B4",X"E0",X"40",X"88",X"44",X"44",X"33",
		X"08",X"4C",X"E8",X"F8",X"F8",X"E8",X"4C",X"08",X"03",X"04",X"04",X"04",X"04",X"04",X"04",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"44",X"00",X"00",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"33",X"11",X"FF",X"77",X"33",X"11",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"F0",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"3C",X"F0",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"87",X"87",X"C3",X"C3",
		X"0F",X"0F",X"0F",X"0F",X"1E",X"1E",X"3C",X"3C",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"C3",X"87",X"87",X"0F",X"0F",X"0F",X"0F",
		X"3C",X"3C",X"1E",X"1E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"C3",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"C3",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",
		X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"00",X"00",X"0E",X"0E",X"0D",X"0F",X"0F",X"0F",X"00",X"40",X"80",X"83",X"87",X"87",X"43",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"4A",X"0F",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",
		X"0F",X"FF",X"0F",X"0D",X"0E",X"0E",X"00",X"00",X"2F",X"53",X"87",X"87",X"83",X"80",X"40",X"00",
		X"0F",X"4A",X"C0",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"30",X"25",X"0F",
		X"00",X"20",X"10",X"1C",X"1E",X"1E",X"AC",X"4F",X"00",X"00",X"07",X"07",X"0B",X"0F",X"FF",X"0F",
		X"0F",X"0F",X"0F",X"03",X"00",X"00",X"00",X"00",X"0F",X"25",X"30",X"00",X"00",X"00",X"00",X"00",
		X"4F",X"2C",X"1E",X"1E",X"1C",X"10",X"20",X"00",X"0F",X"0F",X"0F",X"0B",X"07",X"07",X"00",X"00",
		X"C1",X"2D",X"1F",X"2F",X"2F",X"2F",X"27",X"2F",X"30",X"40",X"01",X"01",X"03",X"03",X"03",X"00",
		X"C0",X"20",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"38",X"4B",X"8F",X"0F",X"0F",X"0F",X"0E",X"0F",
		X"0F",X"0F",X"07",X"07",X"43",X"61",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0E",X"0E",X"2C",X"68",X"0C",X"08",
		X"01",X"03",X"61",X"43",X"07",X"07",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"0C",X"68",X"2C",X"0E",X"0E",X"0F",X"0F",
		X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"2D",X"C1",X"00",X"03",X"03",X"03",X"01",X"81",X"40",X"30",
		X"00",X"0C",X"0C",X"0C",X"08",X"18",X"20",X"C0",X"4F",X"4E",X"4F",X"4F",X"4F",X"8F",X"4B",X"38",
		X"00",X"0F",X"6F",X"4F",X"7F",X"0F",X"7F",X"4F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"EF",X"AF",X"AF",X"0F",X"EF",X"2F",
		X"7F",X"0F",X"7F",X"4F",X"7F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EF",X"0F",X"EF",X"2F",X"EF",X"0F",X"0F",X"00",
		X"00",X"0F",X"6F",X"5F",X"4F",X"0F",X"6F",X"4F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"6F",X"2F",X"EF",X"0F",X"EF",X"AF",
		X"7F",X"0F",X"7F",X"4F",X"7F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"AF",X"0F",X"EF",X"2F",X"EF",X"0F",X"0F",X"00",
		X"00",X"0F",X"0F",X"0F",X"7F",X"0F",X"7F",X"4F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"4F",X"EF",X"0F",X"EF",X"2F",
		X"7F",X"0F",X"7F",X"4F",X"7F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"EF",X"0F",X"EF",X"2F",X"EF",X"0F",X"0F",X"00",
		X"00",X"0F",X"0F",X"0F",X"69",X"4B",X"78",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"0F",X"0F",X"0F",X"E1",X"A5",X"A5",X"0F",
		X"78",X"4B",X"78",X"0F",X"0F",X"0F",X"0F",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"E1",X"2D",X"E1",X"0F",X"0F",X"0F",X"0F",X"00",
		X"0F",X"0F",X"87",X"C3",X"CB",X"E9",X"ED",X"ED",X"0F",X"0F",X"F0",X"FF",X"FF",X"FF",X"F3",X"FF",
		X"ED",X"ED",X"E9",X"CB",X"C3",X"87",X"0F",X"0F",X"FF",X"FF",X"FF",X"FF",X"FF",X"F0",X"0F",X"0F",
		X"FF",X"FF",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"CF",X"9E",X"3C",X"78",X"78",X"78",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"FF",X"FF",X"78",X"78",X"78",X"3C",X"9E",X"CF",X"FF",X"FF",
		X"0F",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"0F",X"08",X"08",X"08",X"1B",X"1B",X"1B",X"1B",
		X"0F",X"01",X"89",X"CD",X"CD",X"CD",X"0D",X"09",X"0F",X"00",X"37",X"37",X"FF",X"F9",X"F7",X"F9",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"0F",X"1B",X"1B",X"1B",X"1B",X"08",X"08",X"08",X"0F",
		X"09",X"0D",X"CD",X"CD",X"CD",X"89",X"01",X"0F",X"FB",X"F5",X"F5",X"FF",X"37",X"37",X"00",X"0F",
		X"0F",X"00",X"EE",X"7F",X"FF",X"EE",X"FF",X"FF",X"0F",X"08",X"3B",X"2A",X"2B",X"3B",X"3B",X"3B",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"81",X"41",X"0F",X"00",X"00",X"00",X"88",X"70",X"88",X"88",
		X"FF",X"FF",X"EE",X"FF",X"FF",X"EE",X"00",X"0F",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"08",X"0F",
		X"41",X"81",X"01",X"01",X"01",X"01",X"01",X"0F",X"88",X"88",X"F0",X"88",X"00",X"00",X"00",X"0F",
		X"0F",X"44",X"E7",X"7F",X"F7",X"7F",X"EE",X"CC",X"0F",X"08",X"18",X"29",X"29",X"29",X"18",X"08",
		X"0F",X"01",X"01",X"81",X"CD",X"CD",X"89",X"89",X"0F",X"00",X"08",X"98",X"FE",X"FF",X"00",X"00",
		X"DD",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"0F",X"08",X"18",X"29",X"29",X"29",X"18",X"08",X"0F",
		X"81",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"88",X"C8",X"C8",X"C8",X"88",X"00",X"00",X"0F",
		X"0F",X"00",X"C0",X"E6",X"EF",X"EF",X"EF",X"EF",X"0F",X"08",X"09",X"09",X"09",X"09",X"09",X"09",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"FC",X"F9",X"F3",X"FF",X"7F",X"3F",X"00",X"0F",X"09",X"09",X"09",X"09",X"09",X"09",X"08",X"0F",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"08",X"8C",X"EC",X"EC",X"EC",X"E8",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"99",X"45",X"02",X"8D",X"0F",X"6E",X"7F",X"3B",X"08",X"08",X"08",X"08",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"89",X"89",X"0F",X"00",X"00",X"00",X"CC",X"37",X"0A",X"05",
		X"8A",X"8D",X"46",X"45",X"33",X"00",X"00",X"0F",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"0F",
		X"4D",X"45",X"4D",X"45",X"89",X"01",X"01",X"0F",X"6E",X"67",X"0A",X"05",X"0A",X"FF",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"BE",X"BE",X"BF",X"C7",X"0F",X"08",X"18",X"18",X"18",X"18",X"18",X"18",
		X"0F",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"00",X"00",X"00",X"00",X"08",X"4C",X"EE",
		X"F7",X"77",X"ED",X"E9",X"8F",X"FF",X"00",X"0F",X"18",X"18",X"19",X"19",X"19",X"19",X"08",X"0F",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"0F",X"EE",X"EE",X"EE",X"EE",X"CC",X"88",X"00",X"0F",
		X"0F",X"00",X"00",X"00",X"80",X"41",X"03",X"17",X"0F",X"4C",X"2A",X"19",X"08",X"08",X"08",X"08",
		X"0F",X"01",X"89",X"CD",X"CD",X"CD",X"CD",X"CD",X"0F",X"00",X"13",X"17",X"3F",X"7F",X"FF",X"DF",
		X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"0F",X"08",X"09",X"0B",X"3B",X"3B",X"19",X"08",X"0F",
		X"89",X"89",X"89",X"01",X"81",X"01",X"01",X"0F",X"EF",X"EF",X"FF",X"FF",X"EE",X"00",X"00",X"0F",
		X"33",X"F3",X"F3",X"F3",X"F3",X"33",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"00",
		X"0F",X"1E",X"3C",X"78",X"F0",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"08",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"FE",X"FE",X"FE",X"FE",X"0F",X"0F",
		X"01",X"01",X"E1",X"EF",X"2F",X"27",X"27",X"27",X"00",X"00",X"F0",X"FF",X"0F",X"08",X"08",X"08",
		X"27",X"2F",X"EF",X"EF",X"E3",X"EB",X"EB",X"EB",X"08",X"0F",X"FF",X"FF",X"F0",X"FF",X"0F",X"0F",
		X"EB",X"EB",X"EB",X"E3",X"EF",X"EF",X"2F",X"27",X"0F",X"0F",X"FF",X"F0",X"FF",X"FF",X"0F",X"08",
		X"27",X"27",X"27",X"2F",X"EF",X"E1",X"01",X"01",X"08",X"08",X"08",X"0F",X"FF",X"F0",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"F0",X"FF",X"3F",X"FF",X"F7",X"F7",X"F7",X"F7",X"F0",X"FF",X"CF",X"FF",
		X"FF",X"3F",X"FF",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"CF",X"FF",X"F0",X"F7",X"F7",X"F7",X"F7",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"55",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"55",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",
		X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"FF",
		X"FF",X"EE",X"FF",X"EE",X"FF",X"EE",X"FF",X"AA",X"77",X"FF",X"77",X"FF",X"77",X"FF",X"77",X"AA",
		X"00",X"11",X"33",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"77",
		X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"AE",X"AE",X"AE",X"00",X"08",X"3D",X"3D",X"3D",X"11",X"00",X"00",
		X"00",X"00",X"8C",X"8F",X"CF",X"CF",X"CF",X"CF",X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",
		X"AE",X"AE",X"AE",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"3D",X"3D",X"3D",X"08",X"00",
		X"CF",X"CF",X"CF",X"CF",X"8F",X"8C",X"00",X"00",X"0C",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"3D",X"3D",X"3D",X"11",X"00",X"00",
		X"00",X"00",X"8E",X"8F",X"CF",X"CF",X"CF",X"CF",X"00",X"00",X"00",X"08",X"4C",X"5F",X"5F",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"3D",X"3D",X"1D",X"18",X"00",
		X"CF",X"CF",X"CF",X"CF",X"8F",X"8E",X"00",X"00",X"5F",X"5F",X"5F",X"4C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"3D",X"3D",X"3D",X"11",X"11",X"11",
		X"00",X"20",X"8E",X"8F",X"8F",X"CF",X"CF",X"CF",X"00",X"00",X"00",X"08",X"4C",X"5F",X"5F",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"3D",X"3D",X"3D",X"08",X"00",
		X"CF",X"CF",X"CF",X"8F",X"8F",X"8E",X"20",X"00",X"5F",X"5F",X"5F",X"4C",X"08",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"08",X"3D",X"3D",X"3D",X"11",X"11",X"11",
		X"00",X"00",X"8B",X"8B",X"8F",X"8F",X"8F",X"8F",X"00",X"80",X"80",X"00",X"6A",X"2F",X"2F",X"2F",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"3D",X"3D",X"3D",X"08",X"00",
		X"8F",X"8F",X"8F",X"8F",X"8B",X"8B",X"00",X"00",X"2F",X"2F",X"2F",X"6A",X"00",X"80",X"80",X"00",
		X"00",X"00",X"00",X"00",X"00",X"4C",X"4C",X"4C",X"00",X"08",X"1D",X"3D",X"3D",X"3D",X"11",X"00",
		X"00",X"00",X"00",X"89",X"CF",X"CF",X"CF",X"CF",X"00",X"20",X"2C",X"0C",X"3D",X"1F",X"1F",X"1F",
		X"4C",X"4C",X"4C",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"3D",X"3D",X"3D",X"1D",X"08",X"00",
		X"CF",X"CF",X"CF",X"CF",X"89",X"00",X"00",X"00",X"1F",X"1F",X"1F",X"3D",X"0C",X"2C",X"20",X"00",
		X"00",X"80",X"80",X"00",X"88",X"AE",X"AE",X"AE",X"00",X"08",X"0C",X"3D",X"3D",X"3D",X"11",X"00",
		X"00",X"00",X"00",X"CC",X"EF",X"EF",X"EF",X"EF",X"00",X"00",X"07",X"07",X"1E",X"0F",X"0F",X"0F",
		X"AE",X"AE",X"AE",X"88",X"00",X"80",X"80",X"00",X"00",X"11",X"3D",X"3D",X"3D",X"0C",X"08",X"00",
		X"EF",X"EF",X"EF",X"EF",X"CC",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"1E",X"07",X"07",X"00",X"00",
		X"00",X"20",X"2C",X"0C",X"C4",X"5F",X"5F",X"5F",X"00",X"00",X"00",X"1D",X"0F",X"0F",X"0F",X"00",
		X"00",X"00",X"00",X"EE",X"FF",X"FF",X"BB",X"33",X"00",X"00",X"01",X"03",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"5F",X"5F",X"C4",X"0C",X"2C",X"20",X"00",X"00",X"07",X"0F",X"0F",X"1D",X"00",X"00",X"00",
		X"33",X"BB",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"03",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"5F",X"D7",X"00",X"0F",X"0F",X"70",X"77",X"77",X"77",X"33",
		X"00",X"00",X"00",X"CF",X"DF",X"DE",X"DE",X"DE",X"00",X"00",X"0C",X"0E",X"8F",X"8F",X"87",X"B4",
		X"5F",X"5F",X"D7",X"5F",X"44",X"00",X"00",X"00",X"00",X"00",X"11",X"3D",X"3D",X"3D",X"0C",X"08",
		X"CF",X"CF",X"CF",X"CF",X"FF",X"B8",X"30",X"00",X"69",X"78",X"7C",X"65",X"10",X"80",X"80",X"00",
		X"08",X"08",X"08",X"08",X"44",X"5F",X"D7",X"5F",X"00",X"01",X"07",X"17",X"17",X"33",X"33",X"11",
		X"00",X"0C",X"0C",X"CC",X"EF",X"EF",X"EF",X"EF",X"F1",X"F3",X"01",X"07",X"0F",X"0F",X"3C",X"69",
		X"5F",X"D7",X"5F",X"44",X"C0",X"C0",X"00",X"00",X"11",X"11",X"33",X"33",X"33",X"30",X"03",X"03",
		X"EF",X"EF",X"EF",X"CD",X"CC",X"80",X"0C",X"0E",X"78",X"7C",X"6D",X"1E",X"2E",X"3E",X"00",X"00",
		X"00",X"00",X"08",X"08",X"C4",X"D7",X"5F",X"D7",X"00",X"00",X"00",X"19",X"1D",X"3D",X"3D",X"2C",
		X"00",X"00",X"DD",X"FE",X"FE",X"FE",X"EF",X"EF",X"00",X"0F",X"8F",X"8F",X"96",X"B4",X"69",X"7C",
		X"D7",X"5F",X"D7",X"C4",X"08",X"08",X"00",X"00",X"00",X"10",X"16",X"16",X"16",X"06",X"04",X"00",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"CC",X"00",X"00",X"7C",X"69",X"3C",X"1E",X"0F",X"FC",X"F8",X"00",
		X"00",X"08",X"0C",X"0C",X"C4",X"5F",X"5F",X"D7",X"00",X"00",X"03",X"07",X"07",X"12",X"11",X"0C",
		X"00",X"00",X"6E",X"7F",X"7F",X"FF",X"FF",X"FF",X"00",X"F1",X"F3",X"0F",X"1E",X"2D",X"7A",X"7A",
		X"D7",X"5F",X"5F",X"C4",X"08",X"08",X"00",X"00",X"3D",X"3D",X"3D",X"19",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"CC",X"00",X"00",X"00",X"7A",X"7A",X"2D",X"1E",X"07",X"E3",X"E3",X"00",
		X"00",X"00",X"00",X"00",X"C4",X"5F",X"5F",X"5F",X"00",X"00",X"00",X"19",X"1D",X"3D",X"3D",X"2C",
		X"00",X"01",X"33",X"F8",X"E9",X"EF",X"EF",X"EF",X"00",X"0C",X"8E",X"8F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"5F",X"5F",X"C4",X"00",X"00",X"00",X"00",X"00",X"33",X"07",X"0F",X"0F",X"0E",X"00",X"00",
		X"EF",X"EF",X"EF",X"EF",X"EF",X"66",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"1E",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"C4",X"5F",X"5F",X"5F",X"00",X"00",X"11",X"33",X"07",X"07",X"03",X"0C",
		X"00",X"00",X"FE",X"EF",X"6F",X"6F",X"6F",X"67",X"00",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"5F",X"5F",X"C4",X"00",X"00",X"00",X"00",X"3D",X"3D",X"3D",X"19",X"00",X"00",X"00",X"00",
		X"EF",X"EF",X"EF",X"EF",X"CC",X"30",X"30",X"00",X"0F",X"0F",X"0F",X"0F",X"07",X"CE",X"C6",X"00",
		X"00",X"00",X"00",X"00",X"C4",X"5F",X"5F",X"5F",X"00",X"00",X"08",X"3D",X"3D",X"3D",X"1D",X"00",
		X"00",X"70",X"71",X"CD",X"EF",X"EF",X"EF",X"EF",X"00",X"8E",X"8F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"5F",X"5F",X"5F",X"C4",X"00",X"00",X"00",X"00",X"00",X"1D",X"3D",X"3D",X"3D",X"08",X"00",X"00",
		X"EF",X"EF",X"EF",X"EF",X"CD",X"71",X"70",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"8F",X"8E",X"00",
		X"00",X"00",X"4C",X"D7",X"5F",X"5F",X"D7",X"5F",X"00",X"00",X"11",X"10",X"10",X"12",X"03",X"33",
		X"00",X"0F",X"8F",X"8F",X"87",X"87",X"0F",X"0F",X"00",X"0E",X"0F",X"1E",X"2D",X"3C",X"78",X"78",
		X"5F",X"44",X"00",X"00",X"00",X"00",X"08",X"0C",X"33",X"33",X"33",X"33",X"33",X"10",X"01",X"01",
		X"EF",X"FF",X"FF",X"FF",X"CC",X"C0",X"0E",X"0F",X"69",X"98",X"EE",X"FF",X"FF",X"70",X"07",X"07",
		X"00",X"44",X"57",X"57",X"57",X"57",X"57",X"57",X"07",X"0F",X"96",X"B4",X"F0",X"3C",X"0F",X"0F",
		X"0C",X"0E",X"C2",X"48",X"E0",X"C0",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"30",X"F8",X"E8",
		X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"33",X"00",
		X"0F",X"0C",X"0C",X"EE",X"FF",X"FF",X"FF",X"77",X"E8",X"00",X"01",X"03",X"83",X"83",X"83",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0C",X"84",X"84",X"00",X"00",X"00",X"01",X"10",X"00",X"11",X"11",
		X"00",X"00",X"0E",X"0D",X"E3",X"EF",X"CF",X"CF",X"00",X"00",X"0E",X"C3",X"C3",X"3C",X"69",X"7C",
		X"84",X"84",X"0C",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"10",X"10",X"01",X"00",X"00",X"00",
		X"CF",X"CF",X"EF",X"E3",X"0D",X"0E",X"00",X"00",X"7C",X"69",X"3C",X"C3",X"C3",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0C",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"31",X"03",
		X"00",X"00",X"21",X"23",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"0F",X"0E",X"EF",X"E9",X"E9",X"0F",
		X"80",X"80",X"84",X"0C",X"08",X"00",X"00",X"00",X"03",X"03",X"03",X"02",X"00",X"00",X"00",X"00",
		X"EF",X"E9",X"E9",X"0F",X"0F",X"07",X"00",X"00",X"3C",X"7A",X"E5",X"D2",X"E1",X"03",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"0C",X"04",X"08",X"00",X"00",X"01",X"03",X"03",X"03",X"02",X"01",
		X"00",X"00",X"B3",X"F7",X"F7",X"FF",X"CF",X"0F",X"00",X"00",X"DC",X"FE",X"FE",X"FF",X"3F",X"0F",
		X"84",X"84",X"0C",X"08",X"00",X"00",X"00",X"00",X"12",X"12",X"03",X"01",X"00",X"00",X"00",X"00",
		X"87",X"B5",X"78",X"5A",X"34",X"07",X"00",X"00",X"1E",X"DA",X"E1",X"A5",X"C2",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"03",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"03",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"0F",X"96",X"B4",X"F0",X"3C",X"0F",X"0F",
		X"88",X"AE",X"AE",X"AE",X"AE",X"AE",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"30",X"F8",X"E8",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"33",X"00",
		X"0F",X"0C",X"0C",X"EE",X"FF",X"FF",X"FF",X"77",X"88",X"00",X"01",X"83",X"C3",X"C3",X"C3",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",
		X"00",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"00",
		X"00",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"30",X"70",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"70",X"30",X"10",X"00",X"00",X"00",X"00",X"00",X"E0",X"F0",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"4A",X"0F",X"00",X"40",X"80",X"83",X"87",X"87",X"43",X"0F",
		X"00",X"00",X"0E",X"0E",X"0D",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0C",X"0F",X"0F",X"0F",
		X"0F",X"4A",X"C0",X"00",X"00",X"00",X"00",X"00",X"2F",X"53",X"87",X"87",X"83",X"80",X"40",X"00",
		X"0F",X"FF",X"0F",X"0D",X"0E",X"0E",X"00",X"00",X"0F",X"0F",X"0F",X"0C",X"00",X"00",X"00",X"00",
		X"00",X"00",X"80",X"00",X"00",X"80",X"84",X"0E",X"00",X"00",X"10",X"60",X"43",X"43",X"03",X"07",
		X"00",X"00",X"07",X"0F",X"0E",X"0F",X"0F",X"0F",X"00",X"10",X"34",X"14",X"0E",X"1E",X"0F",X"0F",
		X"0E",X"84",X"80",X"00",X"00",X"80",X"00",X"00",X"17",X"03",X"43",X"43",X"60",X"10",X"00",X"00",
		X"8F",X"7F",X"0F",X"0E",X"0F",X"07",X"00",X"00",X"0F",X"CF",X"1E",X"0E",X"14",X"34",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"61",X"43",X"07",X"07",X"0F",X"0F",X"08",X"0C",X"68",X"2C",X"0E",X"0E",X"0F",X"0F",
		X"00",X"0C",X"0C",X"0C",X"08",X"08",X"20",X"C0",X"00",X"03",X"03",X"03",X"01",X"01",X"40",X"30",
		X"0F",X"07",X"0F",X"0F",X"0F",X"0F",X"2D",X"C1",X"4F",X"4E",X"4F",X"4F",X"4F",X"8F",X"4B",X"38",
		X"00",X"00",X"00",X"40",X"E0",X"40",X"0C",X"00",X"00",X"00",X"00",X"20",X"70",X"00",X"03",X"00",
		X"00",X"01",X"03",X"61",X"43",X"0F",X"0F",X"0F",X"00",X"08",X"0C",X"68",X"2C",X"0F",X"4F",X"4F",
		X"0C",X"0C",X"0C",X"08",X"40",X"80",X"80",X"00",X"03",X"03",X"03",X"01",X"20",X"10",X"10",X"00",
		X"07",X"0F",X"0F",X"0F",X"0F",X"0F",X"C1",X"00",X"4E",X"4F",X"4F",X"8F",X"8F",X"0F",X"38",X"00",
		X"00",X"00",X"A0",X"70",X"20",X"C0",X"4A",X"0F",X"00",X"00",X"00",X"00",X"08",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"70",X"86",X"0C",X"0F",X"0F",X"0F",
		X"0F",X"4A",X"C0",X"20",X"70",X"A0",X"00",X"00",X"EF",X"1F",X"0F",X"08",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0F",X"CF",X"0F",X"0C",X"86",X"70",X"00",X"00",
		X"00",X"00",X"00",X"0E",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"20",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C3",X"60",X"00",X"00",X"00",
		X"01",X"03",X"07",X"0F",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"10",X"20",X"00",X"00",X"00",X"00",X"60",X"C3",X"00",X"00",X"00",
		X"80",X"C0",X"80",X"40",X"40",X"48",X"48",X"80",X"10",X"30",X"10",X"20",X"20",X"21",X"21",X"10",
		X"01",X"83",X"61",X"43",X"07",X"07",X"0F",X"0F",X"08",X"1C",X"68",X"2C",X"0E",X"0E",X"4F",X"4F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"0F",X"4F",X"4F",X"4F",X"4F",X"4E",X"8E",X"8E",X"8F",
		X"00",X"08",X"08",X"08",X"08",X"08",X"80",X"80",X"00",X"01",X"01",X"01",X"01",X"01",X"10",X"10",
		X"0F",X"0E",X"0C",X"08",X"00",X"80",X"80",X"00",X"0F",X"07",X"03",X"01",X"00",X"10",X"10",X"00",
		X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0C",X"8E",X"86",X"87",X"8F",X"66",X"FF",X"F9",X"F9",X"F9",X"FF",X"67",X"63",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"80",X"FF",X"F9",X"9E",X"FE",X"FF",X"FF",
		X"0F",X"0F",X"0E",X"2F",X"67",X"03",X"00",X"00",X"47",X"CF",X"CB",X"CB",X"E9",X"FF",X"66",X"00",
		X"0F",X"0F",X"1F",X"0F",X"0F",X"07",X"00",X"00",X"7F",X"CF",X"3C",X"3C",X"1F",X"EE",X"FF",X"77",
		X"00",X"00",X"00",X"00",X"8C",X"8E",X"86",X"EE",X"00",X"00",X"01",X"03",X"67",X"FF",X"F9",X"F9",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"80",X"FF",X"9F",X"F8",X"FE",X"7F",
		X"EE",X"FF",X"EE",X"4E",X"CE",X"06",X"00",X"00",X"F9",X"FF",X"EF",X"CB",X"CF",X"67",X"00",X"00",
		X"0F",X"1F",X"2F",X"1F",X"0F",X"0F",X"07",X"00",X"C3",X"F3",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"8C",X"8E",X"86",X"8F",X"66",X"FF",X"F9",X"DB",X"CB",X"CF",X"47",X"03",
		X"44",X"EE",X"EE",X"EF",X"4F",X"4F",X"69",X"69",X"00",X"00",X"80",X"FF",X"F9",X"9E",X"FE",X"FE",
		X"8F",X"0F",X"0F",X"4E",X"CE",X"06",X"00",X"00",X"67",X"FF",X"F9",X"F9",X"F9",X"FF",X"66",X"00",
		X"4F",X"2F",X"2F",X"1F",X"0F",X"0F",X"07",X"00",X"FF",X"7F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",
		X"03",X"47",X"CE",X"0C",X"8E",X"CA",X"C7",X"CF",X"00",X"61",X"47",X"47",X"47",X"43",X"03",X"03",
		X"17",X"69",X"69",X"0F",X"0F",X"0F",X"0F",X"0F",X"88",X"8E",X"0F",X"0F",X"7F",X"FC",X"CF",X"F7",
		X"CF",X"C7",X"CA",X"8E",X"EE",X"FF",X"EF",X"03",X"03",X"03",X"61",X"FF",X"FF",X"FF",X"61",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"1F",X"17",X"F7",X"FC",X"CF",X"7F",X"0F",X"79",X"68",X"88",
		X"8C",X"CE",X"8E",X"0C",X"8E",X"CA",X"C7",X"CF",X"00",X"61",X"FF",X"FF",X"FF",X"61",X"03",X"03",
		X"17",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"4F",X"88",X"68",X"69",X"0F",X"7F",X"CF",X"FC",X"F7",
		X"CF",X"C7",X"CA",X"8E",X"0C",X"8E",X"CE",X"8C",X"13",X"13",X"53",X"47",X"47",X"47",X"61",X"00",
		X"EF",X"EF",X"EF",X"4F",X"4F",X"69",X"69",X"17",X"F7",X"CF",X"FC",X"7F",X"0F",X"0F",X"8E",X"88",
		X"00",X"00",X"00",X"8C",X"8E",X"8E",X"8F",X"8F",X"66",X"FF",X"F9",X"F9",X"F9",X"FF",X"67",X"03",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"69",X"69",X"00",X"80",X"FF",X"9F",X"DB",X"FF",X"FF",X"FF",
		X"0F",X"0F",X"0E",X"2F",X"67",X"03",X"00",X"00",X"47",X"CF",X"CB",X"CB",X"E9",X"FF",X"66",X"00",
		X"4F",X"6F",X"1F",X"0F",X"0F",X"07",X"00",X"00",X"7F",X"0F",X"0F",X"0F",X"0F",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"8C",X"8E",X"8E",X"8F",X"00",X"00",X"01",X"03",X"67",X"FF",X"F9",X"F9",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"80",X"FF",X"D3",X"9F",X"FF",X"FF",
		X"8F",X"0F",X"0F",X"4E",X"CE",X"06",X"00",X"00",X"F9",X"FF",X"EF",X"CB",X"CF",X"67",X"00",X"00",
		X"0F",X"0F",X"0F",X"0F",X"69",X"79",X"07",X"00",X"FF",X"7F",X"0F",X"8F",X"8F",X"8F",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"8C",X"8E",X"8E",X"8F",X"66",X"FF",X"E9",X"CB",X"CB",X"CF",X"47",X"03",
		X"00",X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"FF",X"9F",X"DB",X"FF",X"FF",
		X"8F",X"0F",X"0F",X"4E",X"CE",X"06",X"00",X"00",X"67",X"FF",X"F9",X"F9",X"F9",X"FF",X"66",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"61",X"71",X"FF",X"7F",X"0F",X"0F",X"8F",X"8F",X"8E",X"88",
		X"03",X"47",X"CE",X"0C",X"8E",X"CE",X"CF",X"CF",X"00",X"61",X"FF",X"FF",X"FF",X"61",X"03",X"03",
		X"71",X"69",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"88",X"8E",X"0F",X"0F",X"7F",X"CF",X"ED",X"F7",
		X"CF",X"CF",X"CE",X"8E",X"0C",X"CE",X"47",X"03",X"03",X"03",X"43",X"47",X"47",X"47",X"61",X"00",
		X"0F",X"0F",X"0F",X"69",X"69",X"4F",X"7F",X"07",X"F7",X"CF",X"ED",X"7F",X"0F",X"0F",X"8E",X"08",
		X"8C",X"CE",X"8E",X"0C",X"8E",X"CE",X"CF",X"CF",X"00",X"61",X"47",X"47",X"47",X"43",X"03",X"03",
		X"07",X"7F",X"4F",X"69",X"69",X"0F",X"0F",X"0F",X"08",X"8E",X"0F",X"0F",X"7F",X"ED",X"CF",X"F7",
		X"CF",X"CF",X"CE",X"8E",X"0C",X"8E",X"CE",X"8C",X"03",X"03",X"61",X"FF",X"FF",X"FF",X"61",X"00",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"69",X"71",X"F7",X"ED",X"CF",X"7F",X"0F",X"0F",X"8E",X"88",
		X"00",X"00",X"00",X"44",X"5F",X"D7",X"5F",X"5F",X"07",X"0F",X"78",X"77",X"77",X"FF",X"FF",X"33",
		X"07",X"0F",X"0F",X"8F",X"8F",X"8F",X"8F",X"8F",X"00",X"08",X"0C",X"0F",X"0F",X"3C",X"69",X"78",
		X"D7",X"5F",X"44",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"3D",X"3D",X"3D",X"1D",X"08",X"00",
		X"CF",X"CF",X"CF",X"CD",X"CD",X"88",X"00",X"00",X"78",X"6D",X"18",X"0C",X"CC",X"C0",X"E0",X"C0",
		X"00",X"00",X"22",X"22",X"A2",X"B7",X"F3",X"B7",X"00",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"CC",X"EE",X"EF",X"EF",X"EF",X"00",X"00",X"00",X"00",X"88",X"DC",X"FC",X"FE",
		X"3F",X"7F",X"BF",X"2E",X"2A",X"22",X"00",X"00",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",
		X"FF",X"F1",X"F9",X"DD",X"CD",X"89",X"00",X"00",X"EF",X"CF",X"8F",X"0F",X"0F",X"0E",X"0C",X"00",
		X"00",X"00",X"22",X"22",X"A2",X"B7",X"F3",X"B7",X"00",X"66",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"88",X"CC",X"EE",X"EF",X"EF",X"EB",X"00",X"00",X"C0",X"E0",X"A8",X"DC",X"FC",X"DC",
		X"3F",X"7F",X"BF",X"2E",X"2A",X"22",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",
		X"FB",X"F9",X"F9",X"DD",X"CC",X"88",X"00",X"00",X"EF",X"CF",X"8F",X"8F",X"0F",X"0F",X"06",X"02",
		X"00",X"00",X"00",X"88",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",
		X"00",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"00",X"00",X"11",X"FF",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",X"FF",X"00",X"FF",X"00",X"00",X"FF",X"00",X"00",
		X"E0",X"F0",X"F0",X"F0",X"E0",X"8F",X"2C",X"F8",X"08",X"14",X"3C",X"3C",X"78",X"78",X"F0",X"71",
		X"C0",X"F0",X"F0",X"F0",X"F2",X"F6",X"FE",X"FE",X"07",X"1E",X"3C",X"F0",X"F3",X"F3",X"97",X"92",
		X"F8",X"2C",X"8F",X"E0",X"F0",X"F0",X"F0",X"E0",X"71",X"F0",X"78",X"78",X"3C",X"3C",X"14",X"08",
		X"FE",X"FE",X"F6",X"F2",X"F0",X"F0",X"F0",X"C0",X"D6",X"97",X"F3",X"F3",X"F0",X"3C",X"1E",X"07",
		X"86",X"87",X"C3",X"E1",X"E8",X"8F",X"AC",X"F4",X"10",X"30",X"16",X"07",X"1E",X"78",X"30",X"10",
		X"C0",X"E0",X"F0",X"F0",X"F0",X"F1",X"F3",X"F7",X"70",X"F0",X"F0",X"F0",X"F1",X"F3",X"87",X"C7",
		X"F4",X"AC",X"8F",X"E8",X"E1",X"C3",X"87",X"86",X"10",X"30",X"78",X"1E",X"07",X"16",X"30",X"10",
		X"F7",X"F3",X"F1",X"F0",X"F0",X"F0",X"E0",X"C0",X"C7",X"87",X"F3",X"F1",X"F0",X"F0",X"F0",X"70",
		X"C0",X"68",X"F0",X"F0",X"F0",X"8F",X"2C",X"F8",X"01",X"01",X"03",X"12",X"10",X"30",X"30",X"30",
		X"38",X"3C",X"78",X"F0",X"F0",X"F1",X"F7",X"FF",X"83",X"C3",X"D2",X"F0",X"F3",X"F3",X"97",X"D2",
		X"F8",X"2D",X"8E",X"F0",X"F0",X"F0",X"68",X"C0",X"30",X"30",X"30",X"10",X"12",X"03",X"01",X"01",
		X"FF",X"F7",X"F1",X"F0",X"F0",X"78",X"3C",X"38",X"D6",X"97",X"F3",X"F3",X"F0",X"D2",X"C3",X"83",
		X"00",X"00",X"08",X"C0",X"E4",X"E0",X"C3",X"E1",X"00",X"00",X"03",X"34",X"70",X"70",X"70",X"61",
		X"00",X"02",X"0C",X"E0",X"F0",X"87",X"0F",X"0F",X"00",X"00",X"00",X"20",X"B0",X"F0",X"F0",X"F0",
		X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",X"00",X"30",X"30",X"70",X"70",X"78",X"78",X"34",X"12",
		X"8C",X"84",X"F3",X"B7",X"B4",X"D2",X"F0",X"90",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",
		X"00",X"00",X"08",X"C0",X"E4",X"E0",X"C3",X"E1",X"00",X"01",X"03",X"34",X"70",X"70",X"30",X"30",
		X"00",X"08",X"00",X"C0",X"C3",X"C3",X"C3",X"C3",X"00",X"00",X"00",X"20",X"70",X"F0",X"F0",X"78",
		X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"C0",X"80",X"30",X"30",X"70",X"70",X"78",X"78",X"2C",X"06",
		X"C3",X"87",X"C3",X"F0",X"F0",X"F0",X"F0",X"00",X"3C",X"3C",X"78",X"F0",X"F0",X"D2",X"16",X"34",
		X"00",X"00",X"80",X"C8",X"C0",X"86",X"C2",X"E0",X"00",X"00",X"00",X"00",X"10",X"34",X"38",X"78",
		X"00",X"00",X"00",X"1E",X"96",X"C3",X"C3",X"C3",X"00",X"01",X"50",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"78",X"78",X"78",X"30",X"30",X"10",X"10",X"00",
		X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"F8",X"F0",X"F0",X"F0",X"F0",X"B0",X"07",X"04",
		X"08",X"C0",X"E4",X"E0",X"C3",X"E1",X"F0",X"F0",X"00",X"00",X"00",X"00",X"04",X"09",X"38",X"78",
		X"00",X"00",X"00",X"10",X"1E",X"0F",X"87",X"87",X"00",X"20",X"70",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"F0",X"E0",X"E0",X"E0",X"C0",X"80",X"00",X"00",X"78",X"78",X"70",X"70",X"30",X"30",X"10",X"00",
		X"D2",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"00",X"F8",X"78",X"78",X"34",X"B4",X"30",X"00",X"00",
		X"00",X"08",X"C0",X"E4",X"E0",X"C3",X"E1",X"F0",X"00",X"00",X"00",X"01",X"10",X"30",X"30",X"30",
		X"00",X"00",X"07",X"3C",X"F0",X"F0",X"F0",X"E1",X"00",X"00",X"20",X"70",X"78",X"78",X"3C",X"3C",
		X"78",X"F8",X"E0",X"E0",X"E0",X"40",X"00",X"00",X"30",X"30",X"30",X"30",X"30",X"10",X"00",X"00",
		X"F1",X"F1",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"7C",X"E9",X"E1",X"F0",X"F0",X"F0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"77",X"44",X"77",X"00",X"77",X"44",X"00",X"00",X"EE",X"AA",X"EE",X"00",X"EE",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"00",X"77",X"44",X"77",X"00",X"00",X"00",X"EE",X"00",X"EE",X"22",X"EE",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
